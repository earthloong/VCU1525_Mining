/*
 * Copyright (c) 2017 Sprocket
 *
 * This is free software: you can redistribute it and/or modify
 * it under the terms of the GNU Affero General Public License with
 * additional permissions to the one published by the Free Software
 * Foundation, either version 3 of the License, or (at your option)
 * any later version. For more information see LICENSE.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU Affero General Public License for more details.
 *
 * You should have received a copy of the GNU Affero General Public License
 * along with this program. If not, see <http://www.gnu.org/licenses/>.
 */

module echo512 (
	input clk,
	input [511:0] data,
	output [31:0] hash
);
	
	reg [31:0] h;
	assign hash = h;

	reg [511:0] msg;

	// ROUND 0

	reg  [127:0] i00_00, i00_01, i00_02, i00_03, i00_10, i00_11, i00_12, i00_13, i00_20, i00_21, i00_22, i00_23;
	wire [127:0] o00_00, o00_01, o00_02, o00_03, o00_10, o00_11, o00_12, o00_13, o00_20, o00_21, o00_22, o00_23;

	aes_round r00_00 (clk, i00_00, o00_00);
	aes_round r00_01 (clk, i00_01, o00_01);
	aes_round r00_02 (clk, i00_02, o00_02);
	aes_round r00_03 (clk, i00_03, o00_03);

	aes_round r00_10 (clk, i00_10, o00_10);
	aes_round r00_11 (clk, i00_11, o00_11);
	aes_round r00_12 (clk, i00_12, o00_12);
	aes_round r00_13 (clk, i00_13, o00_13);
	
	echo_mix  r00_20 (clk, i00_20, o00_20);
	echo_mix  r00_21 (clk, i00_21, o00_21);
	echo_mix  r00_22 (clk, i00_22, o00_22);
	echo_mix  r00_23 (clk, i00_23, o00_23);

	always @ ( posedge clk ) begin

		i00_00 <= 128'h00000200000000000000000000000000;
		i00_01 <= 128'h00000200000000000000000000000000;
		i00_02 <= { msg[((2*4)+0)*32 +: 32],	msg[((2*4)+1)*32 +: 32], msg[((2*4)+2)*32 +: 32], msg[((2*4)+3)*32 +: 32] };
		i00_03 <= 128'h00000200000000000000000000000000;

		i00_10 <= { o00_00[127:108], o00_00[107:96] ^ 12'h0200, o00_00[95:0] };
		i00_11 <= { o00_01[127:108], o00_01[107:96] ^ 12'h0205, o00_01[95:0] };
		i00_12 <= { o00_02[127:108], o00_02[107:96] ^ 12'h020A, o00_02[95:0] };
		i00_13 <= { o00_03[127:108], o00_03[107:96] ^ 12'h020F, o00_03[95:0] };

		i00_20 <= { o00_10[127:120], o00_11[127:120], o00_12[127:120], o00_13[127:120], o00_10[119:112], o00_11[119:112], o00_12[119:112], o00_13[119:112], o00_10[111:104], o00_11[111:104], o00_12[111:104], o00_13[111:104], o00_10[103: 96], o00_11[103: 96], o00_12[103: 96], o00_13[103: 96] };
		i00_21 <= { o00_10[ 95: 88], o00_11[ 95: 88], o00_12[ 95: 88], o00_13[ 95: 88], o00_10[ 87: 80], o00_11[ 87: 80], o00_12[ 87: 80], o00_13[ 87: 80], o00_10[ 79: 72], o00_11[ 79: 72], o00_12[ 79: 72], o00_13[ 79: 72],	o00_10[ 71: 64], o00_11[ 71: 64], o00_12[ 71: 64], o00_13[ 71: 64] };
		i00_22 <= { o00_10[ 63: 56], o00_11[ 63: 56], o00_12[ 63: 56], o00_13[ 63: 56], o00_10[ 55: 48], o00_11[ 55: 48], o00_12[ 55: 48], o00_13[ 55: 48], o00_10[ 47: 40], o00_11[ 47: 40], o00_12[ 47: 40], o00_13[ 47: 40], o00_10[ 39: 32], o00_11[ 39: 32], o00_12[ 39: 32], o00_13[ 39: 32] };
		i00_23 <= { o00_10[ 31: 24], o00_11[ 31: 24], o00_12[ 31: 24], o00_13[ 31: 24], o00_10[ 23: 16], o00_11[ 23: 16], o00_12[ 23: 16], o00_13[ 23: 16], o00_10[ 15:  8], o00_11[ 15:  8], o00_12[ 15:  8], o00_13[ 15:  8], o00_10[  7:  0], o00_11[  7:  0], o00_12[  7:  0], o00_13[  7:  0] };
		
	end

	reg  [127:0] i01_00, i01_01, i01_02, i01_03, i01_10, i01_11, i01_12, i01_13, i01_20, i01_21, i01_22, i01_23;
	wire [127:0] o01_00, o01_01, o01_02, o01_03, o01_10, o01_11, o01_12, o01_13, o01_20, o01_21, o01_22, o01_23;

	aes_round r01_00 (clk, i01_00, o01_00);
	aes_round r01_01 (clk, i01_01, o01_01);
	aes_round r01_02 (clk, i01_02, o01_02);
	aes_round r01_03 (clk, i01_03, o01_03);

	aes_round r01_10 (clk, i01_10, o01_10);
	aes_round r01_11 (clk, i01_11, o01_11);
	aes_round r01_12 (clk, i01_12, o01_12);
	aes_round r01_13 (clk, i01_13, o01_13);
	
	echo_mix  r01_20 (clk, i01_20, o01_20);
	echo_mix  r01_21 (clk, i01_21, o01_21);
	echo_mix  r01_22 (clk, i01_22, o01_22);
	echo_mix  r01_23 (clk, i01_23, o01_23);

	always @ ( posedge clk ) begin

		i01_00 <= 128'h00000200000000000000000000000000;
		i01_01 <= { msg[((1*4)+0)*32 +: 32], msg[((1*4)+1)*32 +: 32], msg[((1*4)+2)*32 +: 32], msg[((1*4)+3)*32 +: 32] };
		i01_02 <= 128'h00000000000000000000000002000000;
		i01_03 <= 128'h00000200000000000000000000000000;

		i01_10 <= { o01_00[127:108], o01_00[107:96] ^ 12'h0204, o01_00[95:0] };
		i01_11 <= { o01_01[127:108], o01_01[107:96] ^ 12'h0209, o01_01[95:0] };
		i01_12 <= { o01_02[127:108], o01_02[107:96] ^ 12'h020E, o01_02[95:0] };
		i01_13 <= { o01_03[127:108], o01_03[107:96] ^ 12'h0203, o01_03[95:0] };

		i01_20 <= { o01_10[127:120], o01_11[127:120], o01_12[127:120], o01_13[127:120], o01_10[119:112], o01_11[119:112], o01_12[119:112], o01_13[119:112], o01_10[111:104], o01_11[111:104], o01_12[111:104], o01_13[111:104], o01_10[103: 96], o01_11[103: 96], o01_12[103: 96], o01_13[103: 96] };
		i01_21 <= { o01_10[ 95: 88], o01_11[ 95: 88], o01_12[ 95: 88], o01_13[ 95: 88], o01_10[ 87: 80], o01_11[ 87: 80], o01_12[ 87: 80], o01_13[ 87: 80], o01_10[ 79: 72], o01_11[ 79: 72], o01_12[ 79: 72], o01_13[ 79: 72],	o01_10[ 71: 64], o01_11[ 71: 64], o01_12[ 71: 64], o01_13[ 71: 64] };
		i01_22 <= { o01_10[ 63: 56], o01_11[ 63: 56], o01_12[ 63: 56], o01_13[ 63: 56], o01_10[ 55: 48], o01_11[ 55: 48], o01_12[ 55: 48], o01_13[ 55: 48], o01_10[ 47: 40], o01_11[ 47: 40], o01_12[ 47: 40], o01_13[ 47: 40], o01_10[ 39: 32], o01_11[ 39: 32], o01_12[ 39: 32], o01_13[ 39: 32] };
		i01_23 <= { o01_10[ 31: 24], o01_11[ 31: 24], o01_12[ 31: 24], o01_13[ 31: 24], o01_10[ 23: 16], o01_11[ 23: 16], o01_12[ 23: 16], o01_13[ 23: 16], o01_10[ 15:  8], o01_11[ 15:  8], o01_12[ 15:  8], o01_13[ 15:  8], o01_10[  7:  0], o01_11[  7:  0], o01_12[  7:  0], o01_13[  7:  0] };

	end

	reg  [127:0] i02_00, i02_01, i02_02, i02_03, i02_10, i02_11, i02_12, i02_13, i02_20, i02_21, i02_22, i02_23;
	wire [127:0] o02_00, o02_01, o02_02, o02_03, o02_10, o02_11, o02_12, o02_13, o02_20, o02_21, o02_22, o02_23;

	aes_round r02_00 (clk, i02_00, o02_00);
	aes_round r02_01 (clk, i02_01, o02_01);
	aes_round r02_02 (clk, i02_02, o02_02);
	aes_round r02_03 (clk, i02_03, o02_03);

	aes_round r02_10 (clk, i02_10, o02_10);
	aes_round r02_11 (clk, i02_11, o02_11);
	aes_round r02_12 (clk, i02_12, o02_12);
	aes_round r02_13 (clk, i02_13, o02_13);
	
	echo_mix  r02_20 (clk, i02_20, o02_20);
	echo_mix  r02_21 (clk, i02_21, o02_21);
	echo_mix  r02_22 (clk, i02_22, o02_22);
	echo_mix  r02_23 (clk, i02_23, o02_23);

	always @ ( posedge clk ) begin

		i02_00 <= { msg[((0*4)+0)*32 +: 32], msg[((0*4)+1)*32 +: 32], msg[((0*4)+2)*32 +: 32], msg[((0*4)+3)*32 +: 32] };
		i02_01 <= 128'h00000000000000000000000000000000;
		i02_02 <= 128'h00000200000000000000000000000000;
		i02_03 <= 128'h00000200000000000000000000000000;

		i02_10 <= { o02_00[127:108], o02_00[107:96] ^ 12'h0208, o02_00[95:0] };
		i02_11 <= { o02_01[127:108], o02_01[107:96] ^ 12'h020D, o02_01[95:0] };
		i02_12 <= { o02_02[127:108], o02_02[107:96] ^ 12'h0202, o02_02[95:0] };
		i02_13 <= { o02_03[127:108], o02_03[107:96] ^ 12'h0207, o02_03[95:0] };

		i02_20 <= { o02_10[127:120], o02_11[127:120], o02_12[127:120], o02_13[127:120], o02_10[119:112], o02_11[119:112], o02_12[119:112], o02_13[119:112], o02_10[111:104], o02_11[111:104], o02_12[111:104], o02_13[111:104], o02_10[103: 96], o02_11[103: 96], o02_12[103: 96], o02_13[103: 96] };
		i02_21 <= { o02_10[ 95: 88], o02_11[ 95: 88], o02_12[ 95: 88], o02_13[ 95: 88], o02_10[ 87: 80], o02_11[ 87: 80], o02_12[ 87: 80], o02_13[ 87: 80], o02_10[ 79: 72], o02_11[ 79: 72], o02_12[ 79: 72], o02_13[ 79: 72],	o02_10[ 71: 64], o02_11[ 71: 64], o02_12[ 71: 64], o02_13[ 71: 64] };
		i02_22 <= { o02_10[ 63: 56], o02_11[ 63: 56], o02_12[ 63: 56], o02_13[ 63: 56], o02_10[ 55: 48], o02_11[ 55: 48], o02_12[ 55: 48], o02_13[ 55: 48], o02_10[ 47: 40], o02_11[ 47: 40], o02_12[ 47: 40], o02_13[ 47: 40], o02_10[ 39: 32], o02_11[ 39: 32], o02_12[ 39: 32], o02_13[ 39: 32] };
		i02_23 <= { o02_10[ 31: 24], o02_11[ 31: 24], o02_12[ 31: 24], o02_13[ 31: 24], o02_10[ 23: 16], o02_11[ 23: 16], o02_12[ 23: 16], o02_13[ 23: 16], o02_10[ 15:  8], o02_11[ 15:  8], o02_12[ 15:  8], o02_13[ 15:  8], o02_10[  7:  0], o02_11[  7:  0], o02_12[  7:  0], o02_13[  7:  0] };

	end

	reg  [127:0] i03_00, i03_01, i03_02, i03_03, i03_10, i03_11, i03_12, i03_13, i03_20, i03_21, i03_22, i03_23;
	wire [127:0] o03_00, o03_01, o03_02, o03_03, o03_10, o03_11, o03_12, o03_13, o03_20, o03_21, o03_22, o03_23;

	aes_round r03_00 (clk, i03_00, o03_00);
	aes_round r03_01 (clk, i03_01, o03_01);
	aes_round r03_02 (clk, i03_02, o03_02);
	aes_round r03_03 (clk, i03_03, o03_03);

	aes_round r03_10 (clk, i03_10, o03_10);
	aes_round r03_11 (clk, i03_11, o03_11);
	aes_round r03_12 (clk, i03_12, o03_12);
	aes_round r03_13 (clk, i03_13, o03_13);
	
	echo_mix  r03_20 (clk, i03_20, o03_20);
	echo_mix  r03_21 (clk, i03_21, o03_21);
	echo_mix  r03_22 (clk, i03_22, o03_22);
	echo_mix  r03_23 (clk, i03_23, o03_23);

	always @ ( posedge clk ) begin

		i03_00 <= 128'h00000080000000000000000000000000;
		i03_01 <= 128'h00000200000000000000000000000000;
		i03_02 <= 128'h00000200000000000000000000000000;
		i03_03 <= { msg[((3*4)+0)*32 +: 32], msg[((3*4)+1)*32 +: 32], msg[((3*4)+2)*32 +: 32],	msg[((3*4)+3)*32 +: 32] };

		i03_10 <= { o03_00[127:108], o03_00[107:96] ^ 12'h020C, o03_00[95:0] };
		i03_11 <= { o03_01[127:108], o03_01[107:96] ^ 12'h0201, o03_01[95:0] };
		i03_12 <= { o03_02[127:108], o03_02[107:96] ^ 12'h0206, o03_02[95:0] };
		i03_13 <= { o03_03[127:108], o03_03[107:96] ^ 12'h020B, o03_03[95:0] };

		i03_20 <= { o03_10[127:120], o03_11[127:120], o03_12[127:120], o03_13[127:120], o03_10[119:112], o03_11[119:112], o03_12[119:112], o03_13[119:112], o03_10[111:104], o03_11[111:104], o03_12[111:104], o03_13[111:104], o03_10[103: 96], o03_11[103: 96], o03_12[103: 96], o03_13[103: 96] };
		i03_21 <= { o03_10[ 95: 88], o03_11[ 95: 88], o03_12[ 95: 88], o03_13[ 95: 88], o03_10[ 87: 80], o03_11[ 87: 80], o03_12[ 87: 80], o03_13[ 87: 80], o03_10[ 79: 72], o03_11[ 79: 72], o03_12[ 79: 72], o03_13[ 79: 72],	o03_10[ 71: 64], o03_11[ 71: 64], o03_12[ 71: 64], o03_13[ 71: 64] };
		i03_22 <= { o03_10[ 63: 56], o03_11[ 63: 56], o03_12[ 63: 56], o03_13[ 63: 56], o03_10[ 55: 48], o03_11[ 55: 48], o03_12[ 55: 48], o03_13[ 55: 48], o03_10[ 47: 40], o03_11[ 47: 40], o03_12[ 47: 40], o03_13[ 47: 40], o03_10[ 39: 32], o03_11[ 39: 32], o03_12[ 39: 32], o03_13[ 39: 32] };
		i03_23 <= { o03_10[ 31: 24], o03_11[ 31: 24], o03_12[ 31: 24], o03_13[ 31: 24], o03_10[ 23: 16], o03_11[ 23: 16], o03_12[ 23: 16], o03_13[ 23: 16], o03_10[ 15:  8], o03_11[ 15:  8], o03_12[ 15:  8], o03_13[ 15:  8], o03_10[  7:  0], o03_11[  7:  0], o03_12[  7:  0], o03_13[  7:  0] };

	end

	// ROUND 1

	reg  [127:0] i10_00, i10_01, i10_02, i10_03, i10_10, i10_11, i10_12, i10_13, i10_20, i10_21, i10_22, i10_23;
	wire [127:0] o10_00, o10_01, o10_02, o10_03, o10_10, o10_11, o10_12, o10_13, o10_20, o10_21, o10_22, o10_23;

	aes_round r10_00 (clk, i10_00, o10_00);
	aes_round r10_01 (clk, i10_01, o10_01);
	aes_round r10_02 (clk, i10_02, o10_02);
	aes_round r10_03 (clk, i10_03, o10_03);

	aes_round r10_10 (clk, i10_10, o10_10);
	aes_round r10_11 (clk, i10_11, o10_11);
	aes_round r10_12 (clk, i10_12, o10_12);
	aes_round r10_13 (clk, i10_13, o10_13);
	
	echo_mix  r10_20 (clk, i10_20, o10_20);
	echo_mix  r10_21 (clk, i10_21, o10_21);
	echo_mix  r10_22 (clk, i10_22, o10_22);
	echo_mix  r10_23 (clk, i10_23, o10_23);

	always @ ( posedge clk ) begin

		i10_00 <= { o00_20[127:120], o00_20[95:88], o00_20[63:56], o00_20[31:24], o00_21[127:120], o00_21[95:88], o00_21[63:56], o00_21[31:24], o00_22[127:120], o00_22[95:88], o00_22[63:56], o00_22[31:24], o00_23[127:120], o00_23[95:88], o00_23[63:56], o00_23[31:24] };
		i10_01 <= { o01_20[119:112], o01_20[87:80], o01_20[55:48], o01_20[23:16], o01_21[119:112], o01_21[87:80], o01_21[55:48], o01_21[23:16], o01_22[119:112], o01_22[87:80], o01_22[55:48], o01_22[23:16], o01_23[119:112], o01_23[87:80], o01_23[55:48], o01_23[23:16] };
		i10_02 <= { o02_20[111:104], o02_20[79:72], o02_20[47:40], o02_20[15: 8], o02_21[111:104], o02_21[79:72], o02_21[47:40], o02_21[15: 8], o02_22[111:104], o02_22[79:72], o02_22[47:40], o02_22[15: 8], o02_23[111:104], o02_23[79:72], o02_23[47:40], o02_23[15: 8] };
		i10_03 <= { o03_20[103: 96], o03_20[71:64], o03_20[39:32], o03_20[ 7: 0], o03_21[103: 96], o03_21[71:64], o03_21[39:32], o03_21[ 7: 0], o03_22[103: 96], o03_22[71:64], o03_22[39:32], o03_22[ 7: 0], o03_23[103: 96], o03_23[71:64], o03_23[39:32], o03_23[ 7: 0] }; 

		i10_10 <= { o10_00[127:108], o10_00[107:96] ^ 12'h0210, o10_00[95:0] };
		i10_11 <= { o10_01[127:108], o10_01[107:96] ^ 12'h0215, o10_01[95:0] };
		i10_12 <= { o10_02[127:108], o10_02[107:96] ^ 12'h021A, o10_02[95:0] };
		i10_13 <= { o10_03[127:108], o10_03[107:96] ^ 12'h021F, o10_03[95:0] };

		i10_20 <= { o10_10[127:120], o10_11[127:120], o10_12[127:120], o10_13[127:120], o10_10[119:112], o10_11[119:112], o10_12[119:112], o10_13[119:112], o10_10[111:104], o10_11[111:104], o10_12[111:104], o10_13[111:104], o10_10[103: 96], o10_11[103: 96], o10_12[103: 96], o10_13[103: 96] };
		i10_21 <= { o10_10[ 95: 88], o10_11[ 95: 88], o10_12[ 95: 88], o10_13[ 95: 88], o10_10[ 87: 80], o10_11[ 87: 80], o10_12[ 87: 80], o10_13[ 87: 80], o10_10[ 79: 72], o10_11[ 79: 72], o10_12[ 79: 72], o10_13[ 79: 72],	o10_10[ 71: 64], o10_11[ 71: 64], o10_12[ 71: 64], o10_13[ 71: 64] };
		i10_22 <= { o10_10[ 63: 56], o10_11[ 63: 56], o10_12[ 63: 56], o10_13[ 63: 56], o10_10[ 55: 48], o10_11[ 55: 48], o10_12[ 55: 48], o10_13[ 55: 48], o10_10[ 47: 40], o10_11[ 47: 40], o10_12[ 47: 40], o10_13[ 47: 40], o10_10[ 39: 32], o10_11[ 39: 32], o10_12[ 39: 32], o10_13[ 39: 32] };
		i10_23 <= { o10_10[ 31: 24], o10_11[ 31: 24], o10_12[ 31: 24], o10_13[ 31: 24], o10_10[ 23: 16], o10_11[ 23: 16], o10_12[ 23: 16], o10_13[ 23: 16], o10_10[ 15:  8], o10_11[ 15:  8], o10_12[ 15:  8], o10_13[ 15:  8], o10_10[  7:  0], o10_11[  7:  0], o10_12[  7:  0], o10_13[  7:  0] };
		
	end

	reg  [127:0] i11_00, i11_01, i11_02, i11_03, i11_10, i11_11, i11_12, i11_13, i11_20, i11_21, i11_22, i11_23;
	wire [127:0] o11_00, o11_01, o11_02, o11_03, o11_10, o11_11, o11_12, o11_13, o11_20, o11_21, o11_22, o11_23;

	aes_round r11_00 (clk, i11_00, o11_00);
	aes_round r11_01 (clk, i11_01, o11_01);
	aes_round r11_02 (clk, i11_02, o11_02);
	aes_round r11_03 (clk, i11_03, o11_03);

	aes_round r11_10 (clk, i11_10, o11_10);
	aes_round r11_11 (clk, i11_11, o11_11);
	aes_round r11_12 (clk, i11_12, o11_12);
	aes_round r11_13 (clk, i11_13, o11_13);
	
	echo_mix  r11_20 (clk, i11_20, o11_20);
	echo_mix  r11_21 (clk, i11_21, o11_21);
	echo_mix  r11_22 (clk, i11_22, o11_22);
	echo_mix  r11_23 (clk, i11_23, o11_23);

	always @ ( posedge clk ) begin

		i11_00 <= { o01_20[127:120], o01_20[95:88], o01_20[63:56], o01_20[31:24], o01_21[127:120], o01_21[95:88], o01_21[63:56], o01_21[31:24], o01_22[127:120], o01_22[95:88], o01_22[63:56], o01_22[31:24], o01_23[127:120], o01_23[95:88], o01_23[63:56], o01_23[31:24] };
		i11_01 <= { o02_20[119:112], o02_20[87:80], o02_20[55:48], o02_20[23:16], o02_21[119:112], o02_21[87:80], o02_21[55:48], o02_21[23:16], o02_22[119:112], o02_22[87:80], o02_22[55:48], o02_22[23:16], o02_23[119:112], o02_23[87:80], o02_23[55:48], o02_23[23:16] };
		i11_02 <= { o03_20[111:104], o03_20[79:72], o03_20[47:40], o03_20[15: 8], o03_21[111:104], o03_21[79:72], o03_21[47:40], o03_21[15: 8], o03_22[111:104], o03_22[79:72], o03_22[47:40], o03_22[15: 8], o03_23[111:104], o03_23[79:72], o03_23[47:40], o03_23[15: 8] };
		i11_03 <= { o00_20[103: 96], o00_20[71:64], o00_20[39:32], o00_20[ 7: 0], o00_21[103: 96], o00_21[71:64], o00_21[39:32], o00_21[ 7: 0], o00_22[103: 96], o00_22[71:64], o00_22[39:32], o00_22[ 7: 0], o00_23[103: 96], o00_23[71:64], o00_23[39:32], o00_23[ 7: 0] };

		i11_10 <= { o11_00[127:108], o11_00[107:96] ^ 12'h0214, o11_00[95:0] };
		i11_11 <= { o11_01[127:108], o11_01[107:96] ^ 12'h0219, o11_01[95:0] };
		i11_12 <= { o11_02[127:108], o11_02[107:96] ^ 12'h021E, o11_02[95:0] };
		i11_13 <= { o11_03[127:108], o11_03[107:96] ^ 12'h0213, o11_03[95:0] };

		i11_20 <= { o11_10[127:120], o11_11[127:120], o11_12[127:120], o11_13[127:120], o11_10[119:112], o11_11[119:112], o11_12[119:112], o11_13[119:112], o11_10[111:104], o11_11[111:104], o11_12[111:104], o11_13[111:104], o11_10[103: 96], o11_11[103: 96], o11_12[103: 96], o11_13[103: 96] };
		i11_21 <= { o11_10[ 95: 88], o11_11[ 95: 88], o11_12[ 95: 88], o11_13[ 95: 88], o11_10[ 87: 80], o11_11[ 87: 80], o11_12[ 87: 80], o11_13[ 87: 80], o11_10[ 79: 72], o11_11[ 79: 72], o11_12[ 79: 72], o11_13[ 79: 72],	o11_10[ 71: 64], o11_11[ 71: 64], o11_12[ 71: 64], o11_13[ 71: 64] };
		i11_22 <= { o11_10[ 63: 56], o11_11[ 63: 56], o11_12[ 63: 56], o11_13[ 63: 56], o11_10[ 55: 48], o11_11[ 55: 48], o11_12[ 55: 48], o11_13[ 55: 48], o11_10[ 47: 40], o11_11[ 47: 40], o11_12[ 47: 40], o11_13[ 47: 40], o11_10[ 39: 32], o11_11[ 39: 32], o11_12[ 39: 32], o11_13[ 39: 32] };
		i11_23 <= { o11_10[ 31: 24], o11_11[ 31: 24], o11_12[ 31: 24], o11_13[ 31: 24], o11_10[ 23: 16], o11_11[ 23: 16], o11_12[ 23: 16], o11_13[ 23: 16], o11_10[ 15:  8], o11_11[ 15:  8], o11_12[ 15:  8], o11_13[ 15:  8], o11_10[  7:  0], o11_11[  7:  0], o11_12[  7:  0], o11_13[  7:  0] };

	end

	reg  [127:0] i12_00, i12_01, i12_02, i12_03, i12_10, i12_11, i12_12, i12_13, i12_20, i12_21, i12_22, i12_23;
	wire [127:0] o12_00, o12_01, o12_02, o12_03, o12_10, o12_11, o12_12, o12_13, o12_20, o12_21, o12_22, o12_23;

	aes_round r12_00 (clk, i12_00, o12_00);
	aes_round r12_01 (clk, i12_01, o12_01);
	aes_round r12_02 (clk, i12_02, o12_02);
	aes_round r12_03 (clk, i12_03, o12_03);

	aes_round r12_10 (clk, i12_10, o12_10);
	aes_round r12_11 (clk, i12_11, o12_11);
	aes_round r12_12 (clk, i12_12, o12_12);
	aes_round r12_13 (clk, i12_13, o12_13);
	
	echo_mix  r12_20 (clk, i12_20, o12_20);
	echo_mix  r12_21 (clk, i12_21, o12_21);
	echo_mix  r12_22 (clk, i12_22, o12_22);
	echo_mix  r12_23 (clk, i12_23, o12_23);

	always @ ( posedge clk ) begin

		i12_00 <= { o02_20[127:120], o02_20[95:88], o02_20[63:56], o02_20[31:24], o02_21[127:120], o02_21[95:88], o02_21[63:56], o02_21[31:24], o02_22[127:120], o02_22[95:88], o02_22[63:56], o02_22[31:24], o02_23[127:120], o02_23[95:88], o02_23[63:56], o02_23[31:24] };
		i12_01 <= { o03_20[119:112], o03_20[87:80], o03_20[55:48], o03_20[23:16], o03_21[119:112], o03_21[87:80], o03_21[55:48], o03_21[23:16], o03_22[119:112], o03_22[87:80], o03_22[55:48], o03_22[23:16], o03_23[119:112], o03_23[87:80], o03_23[55:48], o03_23[23:16] };
		i12_02 <= { o00_20[111:104], o00_20[79:72], o00_20[47:40], o00_20[15: 8], o00_21[111:104], o00_21[79:72], o00_21[47:40], o00_21[15: 8], o00_22[111:104], o00_22[79:72], o00_22[47:40], o00_22[15: 8], o00_23[111:104], o00_23[79:72], o00_23[47:40], o00_23[15: 8] };
		i12_03 <= { o01_20[103: 96], o01_20[71:64], o01_20[39:32], o01_20[ 7: 0], o01_21[103: 96], o01_21[71:64], o01_21[39:32], o01_21[ 7: 0], o01_22[103: 96], o01_22[71:64], o01_22[39:32], o01_22[ 7: 0], o01_23[103: 96], o01_23[71:64], o01_23[39:32], o01_23[ 7: 0] }; 

		i12_10 <= { o12_00[127:108], o12_00[107:96] ^ 12'h0218, o12_00[95:0] };
		i12_11 <= { o12_01[127:108], o12_01[107:96] ^ 12'h021D, o12_01[95:0] };
		i12_12 <= { o12_02[127:108], o12_02[107:96] ^ 12'h0212, o12_02[95:0] };
		i12_13 <= { o12_03[127:108], o12_03[107:96] ^ 12'h0217, o12_03[95:0] };

		i12_20 <= { o12_10[127:120], o12_11[127:120], o12_12[127:120], o12_13[127:120], o12_10[119:112], o12_11[119:112], o12_12[119:112], o12_13[119:112], o12_10[111:104], o12_11[111:104], o12_12[111:104], o12_13[111:104], o12_10[103: 96], o12_11[103: 96], o12_12[103: 96], o12_13[103: 96] };
		i12_21 <= { o12_10[ 95: 88], o12_11[ 95: 88], o12_12[ 95: 88], o12_13[ 95: 88], o12_10[ 87: 80], o12_11[ 87: 80], o12_12[ 87: 80], o12_13[ 87: 80], o12_10[ 79: 72], o12_11[ 79: 72], o12_12[ 79: 72], o12_13[ 79: 72],	o12_10[ 71: 64], o12_11[ 71: 64], o12_12[ 71: 64], o12_13[ 71: 64] };
		i12_22 <= { o12_10[ 63: 56], o12_11[ 63: 56], o12_12[ 63: 56], o12_13[ 63: 56], o12_10[ 55: 48], o12_11[ 55: 48], o12_12[ 55: 48], o12_13[ 55: 48], o12_10[ 47: 40], o12_11[ 47: 40], o12_12[ 47: 40], o12_13[ 47: 40], o12_10[ 39: 32], o12_11[ 39: 32], o12_12[ 39: 32], o12_13[ 39: 32] };
		i12_23 <= { o12_10[ 31: 24], o12_11[ 31: 24], o12_12[ 31: 24], o12_13[ 31: 24], o12_10[ 23: 16], o12_11[ 23: 16], o12_12[ 23: 16], o12_13[ 23: 16], o12_10[ 15:  8], o12_11[ 15:  8], o12_12[ 15:  8], o12_13[ 15:  8], o12_10[  7:  0], o12_11[  7:  0], o12_12[  7:  0], o12_13[  7:  0] };

	end

	reg  [127:0] i13_00, i13_01, i13_02, i13_03, i13_10, i13_11, i13_12, i13_13, i13_20, i13_21, i13_22, i13_23;
	wire [127:0] o13_00, o13_01, o13_02, o13_03, o13_10, o13_11, o13_12, o13_13, o13_20, o13_21, o13_22, o13_23;

	aes_round r13_00 (clk, i13_00, o13_00);
	aes_round r13_01 (clk, i13_01, o13_01);
	aes_round r13_02 (clk, i13_02, o13_02);
	aes_round r13_03 (clk, i13_03, o13_03);

	aes_round r13_10 (clk, i13_10, o13_10);
	aes_round r13_11 (clk, i13_11, o13_11);
	aes_round r13_12 (clk, i13_12, o13_12);
	aes_round r13_13 (clk, i13_13, o13_13);
	
	echo_mix  r13_20 (clk, i13_20, o13_20);
	echo_mix  r13_21 (clk, i13_21, o13_21);
	echo_mix  r13_22 (clk, i13_22, o13_22);
	echo_mix  r13_23 (clk, i13_23, o13_23);

	always @ ( posedge clk ) begin

		i13_00 <= { o03_20[127:120], o03_20[95:88], o03_20[63:56], o03_20[31:24], o03_21[127:120], o03_21[95:88], o03_21[63:56], o03_21[31:24], o03_22[127:120], o03_22[95:88], o03_22[63:56], o03_22[31:24], o03_23[127:120], o03_23[95:88], o03_23[63:56], o03_23[31:24] };
		i13_01 <= { o00_20[119:112], o00_20[87:80], o00_20[55:48], o00_20[23:16], o00_21[119:112], o00_21[87:80], o00_21[55:48], o00_21[23:16], o00_22[119:112], o00_22[87:80], o00_22[55:48], o00_22[23:16], o00_23[119:112], o00_23[87:80], o00_23[55:48], o00_23[23:16] };
		i13_02 <= { o01_20[111:104], o01_20[79:72], o01_20[47:40], o01_20[15: 8], o01_21[111:104], o01_21[79:72], o01_21[47:40], o01_21[15: 8], o01_22[111:104], o01_22[79:72], o01_22[47:40], o01_22[15: 8], o01_23[111:104], o01_23[79:72], o01_23[47:40], o01_23[15: 8] };
		i13_03 <= { o02_20[103: 96], o02_20[71:64], o02_20[39:32], o02_20[ 7: 0], o02_21[103: 96], o02_21[71:64], o02_21[39:32], o02_21[ 7: 0], o02_22[103: 96], o02_22[71:64], o02_22[39:32], o02_22[ 7: 0], o02_23[103: 96], o02_23[71:64], o02_23[39:32], o02_23[ 7: 0] }; 

		i13_10 <= { o13_00[127:108], o13_00[107:96] ^ 12'h021C, o13_00[95:0] };
		i13_11 <= { o13_01[127:108], o13_01[107:96] ^ 12'h0211, o13_01[95:0] };
		i13_12 <= { o13_02[127:108], o13_02[107:96] ^ 12'h0216, o13_02[95:0] };
		i13_13 <= { o13_03[127:108], o13_03[107:96] ^ 12'h021B, o13_03[95:0] };

		i13_20 <= { o13_10[127:120], o13_11[127:120], o13_12[127:120], o13_13[127:120], o13_10[119:112], o13_11[119:112], o13_12[119:112], o13_13[119:112], o13_10[111:104], o13_11[111:104], o13_12[111:104], o13_13[111:104], o13_10[103: 96], o13_11[103: 96], o13_12[103: 96], o13_13[103: 96] };
		i13_21 <= { o13_10[ 95: 88], o13_11[ 95: 88], o13_12[ 95: 88], o13_13[ 95: 88], o13_10[ 87: 80], o13_11[ 87: 80], o13_12[ 87: 80], o13_13[ 87: 80], o13_10[ 79: 72], o13_11[ 79: 72], o13_12[ 79: 72], o13_13[ 79: 72],	o13_10[ 71: 64], o13_11[ 71: 64], o13_12[ 71: 64], o13_13[ 71: 64] };
		i13_22 <= { o13_10[ 63: 56], o13_11[ 63: 56], o13_12[ 63: 56], o13_13[ 63: 56], o13_10[ 55: 48], o13_11[ 55: 48], o13_12[ 55: 48], o13_13[ 55: 48], o13_10[ 47: 40], o13_11[ 47: 40], o13_12[ 47: 40], o13_13[ 47: 40], o13_10[ 39: 32], o13_11[ 39: 32], o13_12[ 39: 32], o13_13[ 39: 32] };
		i13_23 <= { o13_10[ 31: 24], o13_11[ 31: 24], o13_12[ 31: 24], o13_13[ 31: 24], o13_10[ 23: 16], o13_11[ 23: 16], o13_12[ 23: 16], o13_13[ 23: 16], o13_10[ 15:  8], o13_11[ 15:  8], o13_12[ 15:  8], o13_13[ 15:  8], o13_10[  7:  0], o13_11[  7:  0], o13_12[  7:  0], o13_13[  7:  0] };

	end

	// ROUND 2

	reg  [127:0] i20_00, i20_01, i20_02, i20_03, i20_10, i20_11, i20_12, i20_13, i20_20, i20_21, i20_22, i20_23;
	wire [127:0] o20_00, o20_01, o20_02, o20_03, o20_10, o20_11, o20_12, o20_13, o20_20, o20_21, o20_22, o20_23;

	aes_round r20_00 (clk, i20_00, o20_00);
	aes_round r20_01 (clk, i20_01, o20_01);
	aes_round r20_02 (clk, i20_02, o20_02);
	aes_round r20_03 (clk, i20_03, o20_03);

	aes_round r20_10 (clk, i20_10, o20_10);
	aes_round r20_11 (clk, i20_11, o20_11);
	aes_round r20_12 (clk, i20_12, o20_12);
	aes_round r20_13 (clk, i20_13, o20_13);
	
	echo_mix  r20_20 (clk, i20_20, o20_20);
	echo_mix  r20_21 (clk, i20_21, o20_21);
	echo_mix  r20_22 (clk, i20_22, o20_22);
	echo_mix  r20_23 (clk, i20_23, o20_23);

	always @ ( posedge clk ) begin

		i20_00 <= { o10_20[127:120], o10_20[95:88], o10_20[63:56], o10_20[31:24], o10_21[127:120], o10_21[95:88], o10_21[63:56], o10_21[31:24], o10_22[127:120], o10_22[95:88], o10_22[63:56], o10_22[31:24], o10_23[127:120], o10_23[95:88], o10_23[63:56], o10_23[31:24] };
		i20_01 <= { o11_20[119:112], o11_20[87:80], o11_20[55:48], o11_20[23:16], o11_21[119:112], o11_21[87:80], o11_21[55:48], o11_21[23:16], o11_22[119:112], o11_22[87:80], o11_22[55:48], o11_22[23:16], o11_23[119:112], o11_23[87:80], o11_23[55:48], o11_23[23:16] };
		i20_02 <= { o12_20[111:104], o12_20[79:72], o12_20[47:40], o12_20[15: 8], o12_21[111:104], o12_21[79:72], o12_21[47:40], o12_21[15: 8], o12_22[111:104], o12_22[79:72], o12_22[47:40], o12_22[15: 8], o12_23[111:104], o12_23[79:72], o12_23[47:40], o12_23[15: 8] };
		i20_03 <= { o13_20[103: 96], o13_20[71:64], o13_20[39:32], o13_20[ 7: 0], o13_21[103: 96], o13_21[71:64], o13_21[39:32], o13_21[ 7: 0], o13_22[103: 96], o13_22[71:64], o13_22[39:32], o13_22[ 7: 0], o13_23[103: 96], o13_23[71:64], o13_23[39:32], o13_23[ 7: 0] }; 

		i20_10 <= { o20_00[127:108], o20_00[107:96] ^ 12'h0220, o20_00[95:0] };
		i20_11 <= { o20_01[127:108], o20_01[107:96] ^ 12'h0225, o20_01[95:0] };
		i20_12 <= { o20_02[127:108], o20_02[107:96] ^ 12'h022A, o20_02[95:0] };
		i20_13 <= { o20_03[127:108], o20_03[107:96] ^ 12'h022F, o20_03[95:0] };

		i20_20 <= { o20_10[127:120], o20_11[127:120], o20_12[127:120], o20_13[127:120], o20_10[119:112], o20_11[119:112], o20_12[119:112], o20_13[119:112], o20_10[111:104], o20_11[111:104], o20_12[111:104], o20_13[111:104], o20_10[103: 96], o20_11[103: 96], o20_12[103: 96], o20_13[103: 96] };
		i20_21 <= { o20_10[ 95: 88], o20_11[ 95: 88], o20_12[ 95: 88], o20_13[ 95: 88], o20_10[ 87: 80], o20_11[ 87: 80], o20_12[ 87: 80], o20_13[ 87: 80], o20_10[ 79: 72], o20_11[ 79: 72], o20_12[ 79: 72], o20_13[ 79: 72],	o20_10[ 71: 64], o20_11[ 71: 64], o20_12[ 71: 64], o20_13[ 71: 64] };
		i20_22 <= { o20_10[ 63: 56], o20_11[ 63: 56], o20_12[ 63: 56], o20_13[ 63: 56], o20_10[ 55: 48], o20_11[ 55: 48], o20_12[ 55: 48], o20_13[ 55: 48], o20_10[ 47: 40], o20_11[ 47: 40], o20_12[ 47: 40], o20_13[ 47: 40], o20_10[ 39: 32], o20_11[ 39: 32], o20_12[ 39: 32], o20_13[ 39: 32] };
		i20_23 <= { o20_10[ 31: 24], o20_11[ 31: 24], o20_12[ 31: 24], o20_13[ 31: 24], o20_10[ 23: 16], o20_11[ 23: 16], o20_12[ 23: 16], o20_13[ 23: 16], o20_10[ 15:  8], o20_11[ 15:  8], o20_12[ 15:  8], o20_13[ 15:  8], o20_10[  7:  0], o20_11[  7:  0], o20_12[  7:  0], o20_13[  7:  0] };
		
	end

	reg  [127:0] i21_00, i21_01, i21_02, i21_03, i21_10, i21_11, i21_12, i21_13, i21_20, i21_21, i21_22, i21_23;
	wire [127:0] o21_00, o21_01, o21_02, o21_03, o21_10, o21_11, o21_12, o21_13, o21_20, o21_21, o21_22, o21_23;

	aes_round r21_00 (clk, i21_00, o21_00);
	aes_round r21_01 (clk, i21_01, o21_01);
	aes_round r21_02 (clk, i21_02, o21_02);
	aes_round r21_03 (clk, i21_03, o21_03);

	aes_round r21_10 (clk, i21_10, o21_10);
	aes_round r21_11 (clk, i21_11, o21_11);
	aes_round r21_12 (clk, i21_12, o21_12);
	aes_round r21_13 (clk, i21_13, o21_13);
	
	echo_mix  r21_20 (clk, i21_20, o21_20);
	echo_mix  r21_21 (clk, i21_21, o21_21);
	echo_mix  r21_22 (clk, i21_22, o21_22);
	echo_mix  r21_23 (clk, i21_23, o21_23);

	always @ ( posedge clk ) begin

		i21_00 <= { o11_20[127:120], o11_20[95:88], o11_20[63:56], o11_20[31:24], o11_21[127:120], o11_21[95:88], o11_21[63:56], o11_21[31:24], o11_22[127:120], o11_22[95:88], o11_22[63:56], o11_22[31:24], o11_23[127:120], o11_23[95:88], o11_23[63:56], o11_23[31:24] };
		i21_01 <= { o12_20[119:112], o12_20[87:80], o12_20[55:48], o12_20[23:16], o12_21[119:112], o12_21[87:80], o12_21[55:48], o12_21[23:16], o12_22[119:112], o12_22[87:80], o12_22[55:48], o12_22[23:16], o12_23[119:112], o12_23[87:80], o12_23[55:48], o12_23[23:16] };
		i21_02 <= { o13_20[111:104], o13_20[79:72], o13_20[47:40], o13_20[15: 8], o13_21[111:104], o13_21[79:72], o13_21[47:40], o13_21[15: 8], o13_22[111:104], o13_22[79:72], o13_22[47:40], o13_22[15: 8], o13_23[111:104], o13_23[79:72], o13_23[47:40], o13_23[15: 8] };
		i21_03 <= { o10_20[103: 96], o10_20[71:64], o10_20[39:32], o10_20[ 7: 0], o10_21[103: 96], o10_21[71:64], o10_21[39:32], o10_21[ 7: 0], o10_22[103: 96], o10_22[71:64], o10_22[39:32], o10_22[ 7: 0], o10_23[103: 96], o10_23[71:64], o10_23[39:32], o10_23[ 7: 0] };

		i21_10 <= { o21_00[127:108], o21_00[107:96] ^ 12'h0224, o21_00[95:0] };
		i21_11 <= { o21_01[127:108], o21_01[107:96] ^ 12'h0229, o21_01[95:0] };
		i21_12 <= { o21_02[127:108], o21_02[107:96] ^ 12'h022E, o21_02[95:0] };
		i21_13 <= { o21_03[127:108], o21_03[107:96] ^ 12'h0223, o21_03[95:0] };

		i21_20 <= { o21_10[127:120], o21_11[127:120], o21_12[127:120], o21_13[127:120], o21_10[119:112], o21_11[119:112], o21_12[119:112], o21_13[119:112], o21_10[111:104], o21_11[111:104], o21_12[111:104], o21_13[111:104], o21_10[103: 96], o21_11[103: 96], o21_12[103: 96], o21_13[103: 96] };
		i21_21 <= { o21_10[ 95: 88], o21_11[ 95: 88], o21_12[ 95: 88], o21_13[ 95: 88], o21_10[ 87: 80], o21_11[ 87: 80], o21_12[ 87: 80], o21_13[ 87: 80], o21_10[ 79: 72], o21_11[ 79: 72], o21_12[ 79: 72], o21_13[ 79: 72],	o21_10[ 71: 64], o21_11[ 71: 64], o21_12[ 71: 64], o21_13[ 71: 64] };
		i21_22 <= { o21_10[ 63: 56], o21_11[ 63: 56], o21_12[ 63: 56], o21_13[ 63: 56], o21_10[ 55: 48], o21_11[ 55: 48], o21_12[ 55: 48], o21_13[ 55: 48], o21_10[ 47: 40], o21_11[ 47: 40], o21_12[ 47: 40], o21_13[ 47: 40], o21_10[ 39: 32], o21_11[ 39: 32], o21_12[ 39: 32], o21_13[ 39: 32] };
		i21_23 <= { o21_10[ 31: 24], o21_11[ 31: 24], o21_12[ 31: 24], o21_13[ 31: 24], o21_10[ 23: 16], o21_11[ 23: 16], o21_12[ 23: 16], o21_13[ 23: 16], o21_10[ 15:  8], o21_11[ 15:  8], o21_12[ 15:  8], o21_13[ 15:  8], o21_10[  7:  0], o21_11[  7:  0], o21_12[  7:  0], o21_13[  7:  0] };

	end

	reg  [127:0] i22_00, i22_01, i22_02, i22_03, i22_10, i22_11, i22_12, i22_13, i22_20, i22_21, i22_22, i22_23;
	wire [127:0] o22_00, o22_01, o22_02, o22_03, o22_10, o22_11, o22_12, o22_13, o22_20, o22_21, o22_22, o22_23;

	aes_round r22_00 (clk, i22_00, o22_00);
	aes_round r22_01 (clk, i22_01, o22_01);
	aes_round r22_02 (clk, i22_02, o22_02);
	aes_round r22_03 (clk, i22_03, o22_03);

	aes_round r22_10 (clk, i22_10, o22_10);
	aes_round r22_11 (clk, i22_11, o22_11);
	aes_round r22_12 (clk, i22_12, o22_12);
	aes_round r22_13 (clk, i22_13, o22_13);
	
	echo_mix  r22_20 (clk, i22_20, o22_20);
	echo_mix  r22_21 (clk, i22_21, o22_21);
	echo_mix  r22_22 (clk, i22_22, o22_22);
	echo_mix  r22_23 (clk, i22_23, o22_23);

	always @ ( posedge clk ) begin

		i22_00 <= { o12_20[127:120], o12_20[95:88], o12_20[63:56], o12_20[31:24], o12_21[127:120], o12_21[95:88], o12_21[63:56], o12_21[31:24], o12_22[127:120], o12_22[95:88], o12_22[63:56], o12_22[31:24], o12_23[127:120], o12_23[95:88], o12_23[63:56], o12_23[31:24] };
		i22_01 <= { o13_20[119:112], o13_20[87:80], o13_20[55:48], o13_20[23:16], o13_21[119:112], o13_21[87:80], o13_21[55:48], o13_21[23:16], o13_22[119:112], o13_22[87:80], o13_22[55:48], o13_22[23:16], o13_23[119:112], o13_23[87:80], o13_23[55:48], o13_23[23:16] };
		i22_02 <= { o10_20[111:104], o10_20[79:72], o10_20[47:40], o10_20[15: 8], o10_21[111:104], o10_21[79:72], o10_21[47:40], o10_21[15: 8], o10_22[111:104], o10_22[79:72], o10_22[47:40], o10_22[15: 8], o10_23[111:104], o10_23[79:72], o10_23[47:40], o10_23[15: 8] };
		i22_03 <= { o11_20[103: 96], o11_20[71:64], o11_20[39:32], o11_20[ 7: 0], o11_21[103: 96], o11_21[71:64], o11_21[39:32], o11_21[ 7: 0], o11_22[103: 96], o11_22[71:64], o11_22[39:32], o11_22[ 7: 0], o11_23[103: 96], o11_23[71:64], o11_23[39:32], o11_23[ 7: 0] }; 

		i22_10 <= { o22_00[127:108], o22_00[107:96] ^ 12'h0228, o22_00[95:0] };
		i22_11 <= { o22_01[127:108], o22_01[107:96] ^ 12'h022D, o22_01[95:0] };
		i22_12 <= { o22_02[127:108], o22_02[107:96] ^ 12'h0222, o22_02[95:0] };
		i22_13 <= { o22_03[127:108], o22_03[107:96] ^ 12'h0227, o22_03[95:0] };

		i22_20 <= { o22_10[127:120], o22_11[127:120], o22_12[127:120], o22_13[127:120], o22_10[119:112], o22_11[119:112], o22_12[119:112], o22_13[119:112], o22_10[111:104], o22_11[111:104], o22_12[111:104], o22_13[111:104], o22_10[103: 96], o22_11[103: 96], o22_12[103: 96], o22_13[103: 96] };
		i22_21 <= { o22_10[ 95: 88], o22_11[ 95: 88], o22_12[ 95: 88], o22_13[ 95: 88], o22_10[ 87: 80], o22_11[ 87: 80], o22_12[ 87: 80], o22_13[ 87: 80], o22_10[ 79: 72], o22_11[ 79: 72], o22_12[ 79: 72], o22_13[ 79: 72],	o22_10[ 71: 64], o22_11[ 71: 64], o22_12[ 71: 64], o22_13[ 71: 64] };
		i22_22 <= { o22_10[ 63: 56], o22_11[ 63: 56], o22_12[ 63: 56], o22_13[ 63: 56], o22_10[ 55: 48], o22_11[ 55: 48], o22_12[ 55: 48], o22_13[ 55: 48], o22_10[ 47: 40], o22_11[ 47: 40], o22_12[ 47: 40], o22_13[ 47: 40], o22_10[ 39: 32], o22_11[ 39: 32], o22_12[ 39: 32], o22_13[ 39: 32] };
		i22_23 <= { o22_10[ 31: 24], o22_11[ 31: 24], o22_12[ 31: 24], o22_13[ 31: 24], o22_10[ 23: 16], o22_11[ 23: 16], o22_12[ 23: 16], o22_13[ 23: 16], o22_10[ 15:  8], o22_11[ 15:  8], o22_12[ 15:  8], o22_13[ 15:  8], o22_10[  7:  0], o22_11[  7:  0], o22_12[  7:  0], o22_13[  7:  0] };

	end

	reg  [127:0] i23_00, i23_01, i23_02, i23_03, i23_10, i23_11, i23_12, i23_13, i23_20, i23_21, i23_22, i23_23;
	wire [127:0] o23_00, o23_01, o23_02, o23_03, o23_10, o23_11, o23_12, o23_13, o23_20, o23_21, o23_22, o23_23;

	aes_round r23_00 (clk, i23_00, o23_00);
	aes_round r23_01 (clk, i23_01, o23_01);
	aes_round r23_02 (clk, i23_02, o23_02);
	aes_round r23_03 (clk, i23_03, o23_03);

	aes_round r23_10 (clk, i23_10, o23_10);
	aes_round r23_11 (clk, i23_11, o23_11);
	aes_round r23_12 (clk, i23_12, o23_12);
	aes_round r23_13 (clk, i23_13, o23_13);
	
	echo_mix  r23_20 (clk, i23_20, o23_20);
	echo_mix  r23_21 (clk, i23_21, o23_21);
	echo_mix  r23_22 (clk, i23_22, o23_22);
	echo_mix  r23_23 (clk, i23_23, o23_23);

	always @ ( posedge clk ) begin

		i23_00 <= { o13_20[127:120], o13_20[95:88], o13_20[63:56], o13_20[31:24], o13_21[127:120], o13_21[95:88], o13_21[63:56], o13_21[31:24], o13_22[127:120], o13_22[95:88], o13_22[63:56], o13_22[31:24], o13_23[127:120], o13_23[95:88], o13_23[63:56], o13_23[31:24] };
		i23_01 <= { o10_20[119:112], o10_20[87:80], o10_20[55:48], o10_20[23:16], o10_21[119:112], o10_21[87:80], o10_21[55:48], o10_21[23:16], o10_22[119:112], o10_22[87:80], o10_22[55:48], o10_22[23:16], o10_23[119:112], o10_23[87:80], o10_23[55:48], o10_23[23:16] };
		i23_02 <= { o11_20[111:104], o11_20[79:72], o11_20[47:40], o11_20[15: 8], o11_21[111:104], o11_21[79:72], o11_21[47:40], o11_21[15: 8], o11_22[111:104], o11_22[79:72], o11_22[47:40], o11_22[15: 8], o11_23[111:104], o11_23[79:72], o11_23[47:40], o11_23[15: 8] };
		i23_03 <= { o12_20[103: 96], o12_20[71:64], o12_20[39:32], o12_20[ 7: 0], o12_21[103: 96], o12_21[71:64], o12_21[39:32], o12_21[ 7: 0], o12_22[103: 96], o12_22[71:64], o12_22[39:32], o12_22[ 7: 0], o12_23[103: 96], o12_23[71:64], o12_23[39:32], o12_23[ 7: 0] }; 

		i23_10 <= { o23_00[127:108], o23_00[107:96] ^ 12'h022C, o23_00[95:0] };
		i23_11 <= { o23_01[127:108], o23_01[107:96] ^ 12'h0221, o23_01[95:0] };
		i23_12 <= { o23_02[127:108], o23_02[107:96] ^ 12'h0226, o23_02[95:0] };
		i23_13 <= { o23_03[127:108], o23_03[107:96] ^ 12'h022B, o23_03[95:0] };

		i23_20 <= { o23_10[127:120], o23_11[127:120], o23_12[127:120], o23_13[127:120], o23_10[119:112], o23_11[119:112], o23_12[119:112], o23_13[119:112], o23_10[111:104], o23_11[111:104], o23_12[111:104], o23_13[111:104], o23_10[103: 96], o23_11[103: 96], o23_12[103: 96], o23_13[103: 96] };
		i23_21 <= { o23_10[ 95: 88], o23_11[ 95: 88], o23_12[ 95: 88], o23_13[ 95: 88], o23_10[ 87: 80], o23_11[ 87: 80], o23_12[ 87: 80], o23_13[ 87: 80], o23_10[ 79: 72], o23_11[ 79: 72], o23_12[ 79: 72], o23_13[ 79: 72],	o23_10[ 71: 64], o23_11[ 71: 64], o23_12[ 71: 64], o23_13[ 71: 64] };
		i23_22 <= { o23_10[ 63: 56], o23_11[ 63: 56], o23_12[ 63: 56], o23_13[ 63: 56], o23_10[ 55: 48], o23_11[ 55: 48], o23_12[ 55: 48], o23_13[ 55: 48], o23_10[ 47: 40], o23_11[ 47: 40], o23_12[ 47: 40], o23_13[ 47: 40], o23_10[ 39: 32], o23_11[ 39: 32], o23_12[ 39: 32], o23_13[ 39: 32] };
		i23_23 <= { o23_10[ 31: 24], o23_11[ 31: 24], o23_12[ 31: 24], o23_13[ 31: 24], o23_10[ 23: 16], o23_11[ 23: 16], o23_12[ 23: 16], o23_13[ 23: 16], o23_10[ 15:  8], o23_11[ 15:  8], o23_12[ 15:  8], o23_13[ 15:  8], o23_10[  7:  0], o23_11[  7:  0], o23_12[  7:  0], o23_13[  7:  0] };

	end

	// ROUND 3

	reg  [127:0] i30_00, i30_01, i30_02, i30_03, i30_10, i30_11, i30_12, i30_13, i30_20, i30_21, i30_22, i30_23;
	wire [127:0] o30_00, o30_01, o30_02, o30_03, o30_10, o30_11, o30_12, o30_13, o30_20, o30_21, o30_22, o30_23;

	aes_round r30_00 (clk, i30_00, o30_00);
	aes_round r30_01 (clk, i30_01, o30_01);
	aes_round r30_02 (clk, i30_02, o30_02);
	aes_round r30_03 (clk, i30_03, o30_03);

	aes_round r30_10 (clk, i30_10, o30_10);
	aes_round r30_11 (clk, i30_11, o30_11);
	aes_round r30_12 (clk, i30_12, o30_12);
	aes_round r30_13 (clk, i30_13, o30_13);
	
	echo_mix  r30_20 (clk, i30_20, o30_20);
	echo_mix  r30_21 (clk, i30_21, o30_21);
	echo_mix  r30_22 (clk, i30_22, o30_22);
	echo_mix  r30_23 (clk, i30_23, o30_23);

	always @ ( posedge clk ) begin

		i30_00 <= { o20_20[127:120], o20_20[95:88], o20_20[63:56], o20_20[31:24], o20_21[127:120], o20_21[95:88], o20_21[63:56], o20_21[31:24], o20_22[127:120], o20_22[95:88], o20_22[63:56], o20_22[31:24], o20_23[127:120], o20_23[95:88], o20_23[63:56], o20_23[31:24] };
		i30_01 <= { o21_20[119:112], o21_20[87:80], o21_20[55:48], o21_20[23:16], o21_21[119:112], o21_21[87:80], o21_21[55:48], o21_21[23:16], o21_22[119:112], o21_22[87:80], o21_22[55:48], o21_22[23:16], o21_23[119:112], o21_23[87:80], o21_23[55:48], o21_23[23:16] };
		i30_02 <= { o22_20[111:104], o22_20[79:72], o22_20[47:40], o22_20[15: 8], o22_21[111:104], o22_21[79:72], o22_21[47:40], o22_21[15: 8], o22_22[111:104], o22_22[79:72], o22_22[47:40], o22_22[15: 8], o22_23[111:104], o22_23[79:72], o22_23[47:40], o22_23[15: 8] };
		i30_03 <= { o23_20[103: 96], o23_20[71:64], o23_20[39:32], o23_20[ 7: 0], o23_21[103: 96], o23_21[71:64], o23_21[39:32], o23_21[ 7: 0], o23_22[103: 96], o23_22[71:64], o23_22[39:32], o23_22[ 7: 0], o23_23[103: 96], o23_23[71:64], o23_23[39:32], o23_23[ 7: 0] }; 

		i30_10 <= { o30_00[127:108], o30_00[107:96] ^ 12'h0230, o30_00[95:0] };
		i30_11 <= { o30_01[127:108], o30_01[107:96] ^ 12'h0235, o30_01[95:0] };
		i30_12 <= { o30_02[127:108], o30_02[107:96] ^ 12'h023A, o30_02[95:0] };
		i30_13 <= { o30_03[127:108], o30_03[107:96] ^ 12'h023F, o30_03[95:0] };

		i30_20 <= { o30_10[127:120], o30_11[127:120], o30_12[127:120], o30_13[127:120], o30_10[119:112], o30_11[119:112], o30_12[119:112], o30_13[119:112], o30_10[111:104], o30_11[111:104], o30_12[111:104], o30_13[111:104], o30_10[103: 96], o30_11[103: 96], o30_12[103: 96], o30_13[103: 96] };
		i30_21 <= { o30_10[ 95: 88], o30_11[ 95: 88], o30_12[ 95: 88], o30_13[ 95: 88], o30_10[ 87: 80], o30_11[ 87: 80], o30_12[ 87: 80], o30_13[ 87: 80], o30_10[ 79: 72], o30_11[ 79: 72], o30_12[ 79: 72], o30_13[ 79: 72],	o30_10[ 71: 64], o30_11[ 71: 64], o30_12[ 71: 64], o30_13[ 71: 64] };
		i30_22 <= { o30_10[ 63: 56], o30_11[ 63: 56], o30_12[ 63: 56], o30_13[ 63: 56], o30_10[ 55: 48], o30_11[ 55: 48], o30_12[ 55: 48], o30_13[ 55: 48], o30_10[ 47: 40], o30_11[ 47: 40], o30_12[ 47: 40], o30_13[ 47: 40], o30_10[ 39: 32], o30_11[ 39: 32], o30_12[ 39: 32], o30_13[ 39: 32] };
		i30_23 <= { o30_10[ 31: 24], o30_11[ 31: 24], o30_12[ 31: 24], o30_13[ 31: 24], o30_10[ 23: 16], o30_11[ 23: 16], o30_12[ 23: 16], o30_13[ 23: 16], o30_10[ 15:  8], o30_11[ 15:  8], o30_12[ 15:  8], o30_13[ 15:  8], o30_10[  7:  0], o30_11[  7:  0], o30_12[  7:  0], o30_13[  7:  0] };
		
	end

	reg  [127:0] i31_00, i31_01, i31_02, i31_03, i31_10, i31_11, i31_12, i31_13, i31_20, i31_21, i31_22, i31_23;
	wire [127:0] o31_00, o31_01, o31_02, o31_03, o31_10, o31_11, o31_12, o31_13, o31_20, o31_21, o31_22, o31_23;

	aes_round r31_00 (clk, i31_00, o31_00);
	aes_round r31_01 (clk, i31_01, o31_01);
	aes_round r31_02 (clk, i31_02, o31_02);
	aes_round r31_03 (clk, i31_03, o31_03);

	aes_round r31_10 (clk, i31_10, o31_10);
	aes_round r31_11 (clk, i31_11, o31_11);
	aes_round r31_12 (clk, i31_12, o31_12);
	aes_round r31_13 (clk, i31_13, o31_13);
	
	echo_mix  r31_20 (clk, i31_20, o31_20);
	echo_mix  r31_21 (clk, i31_21, o31_21);
	echo_mix  r31_22 (clk, i31_22, o31_22);
	echo_mix  r31_23 (clk, i31_23, o31_23);

	always @ ( posedge clk ) begin

		i31_00 <= { o21_20[127:120], o21_20[95:88], o21_20[63:56], o21_20[31:24], o21_21[127:120], o21_21[95:88], o21_21[63:56], o21_21[31:24], o21_22[127:120], o21_22[95:88], o21_22[63:56], o21_22[31:24], o21_23[127:120], o21_23[95:88], o21_23[63:56], o21_23[31:24] };
		i31_01 <= { o22_20[119:112], o22_20[87:80], o22_20[55:48], o22_20[23:16], o22_21[119:112], o22_21[87:80], o22_21[55:48], o22_21[23:16], o22_22[119:112], o22_22[87:80], o22_22[55:48], o22_22[23:16], o22_23[119:112], o22_23[87:80], o22_23[55:48], o22_23[23:16] };
		i31_02 <= { o23_20[111:104], o23_20[79:72], o23_20[47:40], o23_20[15: 8], o23_21[111:104], o23_21[79:72], o23_21[47:40], o23_21[15: 8], o23_22[111:104], o23_22[79:72], o23_22[47:40], o23_22[15: 8], o23_23[111:104], o23_23[79:72], o23_23[47:40], o23_23[15: 8] };
		i31_03 <= { o20_20[103: 96], o20_20[71:64], o20_20[39:32], o20_20[ 7: 0], o20_21[103: 96], o20_21[71:64], o20_21[39:32], o20_21[ 7: 0], o20_22[103: 96], o20_22[71:64], o20_22[39:32], o20_22[ 7: 0], o20_23[103: 96], o20_23[71:64], o20_23[39:32], o20_23[ 7: 0] };

		i31_10 <= { o31_00[127:108], o31_00[107:96] ^ 12'h0234, o31_00[95:0] };
		i31_11 <= { o31_01[127:108], o31_01[107:96] ^ 12'h0239, o31_01[95:0] };
		i31_12 <= { o31_02[127:108], o31_02[107:96] ^ 12'h023E, o31_02[95:0] };
		i31_13 <= { o31_03[127:108], o31_03[107:96] ^ 12'h0233, o31_03[95:0] };

		i31_20 <= { o31_10[127:120], o31_11[127:120], o31_12[127:120], o31_13[127:120], o31_10[119:112], o31_11[119:112], o31_12[119:112], o31_13[119:112], o31_10[111:104], o31_11[111:104], o31_12[111:104], o31_13[111:104], o31_10[103: 96], o31_11[103: 96], o31_12[103: 96], o31_13[103: 96] };
		i31_21 <= { o31_10[ 95: 88], o31_11[ 95: 88], o31_12[ 95: 88], o31_13[ 95: 88], o31_10[ 87: 80], o31_11[ 87: 80], o31_12[ 87: 80], o31_13[ 87: 80], o31_10[ 79: 72], o31_11[ 79: 72], o31_12[ 79: 72], o31_13[ 79: 72],	o31_10[ 71: 64], o31_11[ 71: 64], o31_12[ 71: 64], o31_13[ 71: 64] };
		i31_22 <= { o31_10[ 63: 56], o31_11[ 63: 56], o31_12[ 63: 56], o31_13[ 63: 56], o31_10[ 55: 48], o31_11[ 55: 48], o31_12[ 55: 48], o31_13[ 55: 48], o31_10[ 47: 40], o31_11[ 47: 40], o31_12[ 47: 40], o31_13[ 47: 40], o31_10[ 39: 32], o31_11[ 39: 32], o31_12[ 39: 32], o31_13[ 39: 32] };
		i31_23 <= { o31_10[ 31: 24], o31_11[ 31: 24], o31_12[ 31: 24], o31_13[ 31: 24], o31_10[ 23: 16], o31_11[ 23: 16], o31_12[ 23: 16], o31_13[ 23: 16], o31_10[ 15:  8], o31_11[ 15:  8], o31_12[ 15:  8], o31_13[ 15:  8], o31_10[  7:  0], o31_11[  7:  0], o31_12[  7:  0], o31_13[  7:  0] };

	end

	reg  [127:0] i32_00, i32_01, i32_02, i32_03, i32_10, i32_11, i32_12, i32_13, i32_20, i32_21, i32_22, i32_23;
	wire [127:0] o32_00, o32_01, o32_02, o32_03, o32_10, o32_11, o32_12, o32_13, o32_20, o32_21, o32_22, o32_23;

	aes_round r32_00 (clk, i32_00, o32_00);
	aes_round r32_01 (clk, i32_01, o32_01);
	aes_round r32_02 (clk, i32_02, o32_02);
	aes_round r32_03 (clk, i32_03, o32_03);

	aes_round r32_10 (clk, i32_10, o32_10);
	aes_round r32_11 (clk, i32_11, o32_11);
	aes_round r32_12 (clk, i32_12, o32_12);
	aes_round r32_13 (clk, i32_13, o32_13);
	
	echo_mix  r32_20 (clk, i32_20, o32_20);
	echo_mix  r32_21 (clk, i32_21, o32_21);
	echo_mix  r32_22 (clk, i32_22, o32_22);
	echo_mix  r32_23 (clk, i32_23, o32_23);

	always @ ( posedge clk ) begin

		i32_00 <= { o22_20[127:120], o22_20[95:88], o22_20[63:56], o22_20[31:24], o22_21[127:120], o22_21[95:88], o22_21[63:56], o22_21[31:24], o22_22[127:120], o22_22[95:88], o22_22[63:56], o22_22[31:24], o22_23[127:120], o22_23[95:88], o22_23[63:56], o22_23[31:24] };
		i32_01 <= { o23_20[119:112], o23_20[87:80], o23_20[55:48], o23_20[23:16], o23_21[119:112], o23_21[87:80], o23_21[55:48], o23_21[23:16], o23_22[119:112], o23_22[87:80], o23_22[55:48], o23_22[23:16], o23_23[119:112], o23_23[87:80], o23_23[55:48], o23_23[23:16] };
		i32_02 <= { o20_20[111:104], o20_20[79:72], o20_20[47:40], o20_20[15: 8], o20_21[111:104], o20_21[79:72], o20_21[47:40], o20_21[15: 8], o20_22[111:104], o20_22[79:72], o20_22[47:40], o20_22[15: 8], o20_23[111:104], o20_23[79:72], o20_23[47:40], o20_23[15: 8] };
		i32_03 <= { o21_20[103: 96], o21_20[71:64], o21_20[39:32], o21_20[ 7: 0], o21_21[103: 96], o21_21[71:64], o21_21[39:32], o21_21[ 7: 0], o21_22[103: 96], o21_22[71:64], o21_22[39:32], o21_22[ 7: 0], o21_23[103: 96], o21_23[71:64], o21_23[39:32], o21_23[ 7: 0] }; 

		i32_10 <= { o32_00[127:108], o32_00[107:96] ^ 12'h0238, o32_00[95:0] };
		i32_11 <= { o32_01[127:108], o32_01[107:96] ^ 12'h023D, o32_01[95:0] };
		i32_12 <= { o32_02[127:108], o32_02[107:96] ^ 12'h0232, o32_02[95:0] };
		i32_13 <= { o32_03[127:108], o32_03[107:96] ^ 12'h0237, o32_03[95:0] };

		i32_20 <= { o32_10[127:120], o32_11[127:120], o32_12[127:120], o32_13[127:120], o32_10[119:112], o32_11[119:112], o32_12[119:112], o32_13[119:112], o32_10[111:104], o32_11[111:104], o32_12[111:104], o32_13[111:104], o32_10[103: 96], o32_11[103: 96], o32_12[103: 96], o32_13[103: 96] };
		i32_21 <= { o32_10[ 95: 88], o32_11[ 95: 88], o32_12[ 95: 88], o32_13[ 95: 88], o32_10[ 87: 80], o32_11[ 87: 80], o32_12[ 87: 80], o32_13[ 87: 80], o32_10[ 79: 72], o32_11[ 79: 72], o32_12[ 79: 72], o32_13[ 79: 72],	o32_10[ 71: 64], o32_11[ 71: 64], o32_12[ 71: 64], o32_13[ 71: 64] };
		i32_22 <= { o32_10[ 63: 56], o32_11[ 63: 56], o32_12[ 63: 56], o32_13[ 63: 56], o32_10[ 55: 48], o32_11[ 55: 48], o32_12[ 55: 48], o32_13[ 55: 48], o32_10[ 47: 40], o32_11[ 47: 40], o32_12[ 47: 40], o32_13[ 47: 40], o32_10[ 39: 32], o32_11[ 39: 32], o32_12[ 39: 32], o32_13[ 39: 32] };
		i32_23 <= { o32_10[ 31: 24], o32_11[ 31: 24], o32_12[ 31: 24], o32_13[ 31: 24], o32_10[ 23: 16], o32_11[ 23: 16], o32_12[ 23: 16], o32_13[ 23: 16], o32_10[ 15:  8], o32_11[ 15:  8], o32_12[ 15:  8], o32_13[ 15:  8], o32_10[  7:  0], o32_11[  7:  0], o32_12[  7:  0], o32_13[  7:  0] };

	end

	reg  [127:0] i33_00, i33_01, i33_02, i33_03, i33_10, i33_11, i33_12, i33_13, i33_20, i33_21, i33_22, i33_23;
	wire [127:0] o33_00, o33_01, o33_02, o33_03, o33_10, o33_11, o33_12, o33_13, o33_20, o33_21, o33_22, o33_23;

	aes_round r33_00 (clk, i33_00, o33_00);
	aes_round r33_01 (clk, i33_01, o33_01);
	aes_round r33_02 (clk, i33_02, o33_02);
	aes_round r33_03 (clk, i33_03, o33_03);

	aes_round r33_10 (clk, i33_10, o33_10);
	aes_round r33_11 (clk, i33_11, o33_11);
	aes_round r33_12 (clk, i33_12, o33_12);
	aes_round r33_13 (clk, i33_13, o33_13);
	
	echo_mix  r33_20 (clk, i33_20, o33_20);
	echo_mix  r33_21 (clk, i33_21, o33_21);
	echo_mix  r33_22 (clk, i33_22, o33_22);
	echo_mix  r33_23 (clk, i33_23, o33_23);

	always @ ( posedge clk ) begin

		i33_00 <= { o23_20[127:120], o23_20[95:88], o23_20[63:56], o23_20[31:24], o23_21[127:120], o23_21[95:88], o23_21[63:56], o23_21[31:24], o23_22[127:120], o23_22[95:88], o23_22[63:56], o23_22[31:24], o23_23[127:120], o23_23[95:88], o23_23[63:56], o23_23[31:24] };
		i33_01 <= { o20_20[119:112], o20_20[87:80], o20_20[55:48], o20_20[23:16], o20_21[119:112], o20_21[87:80], o20_21[55:48], o20_21[23:16], o20_22[119:112], o20_22[87:80], o20_22[55:48], o20_22[23:16], o20_23[119:112], o20_23[87:80], o20_23[55:48], o20_23[23:16] };
		i33_02 <= { o21_20[111:104], o21_20[79:72], o21_20[47:40], o21_20[15: 8], o21_21[111:104], o21_21[79:72], o21_21[47:40], o21_21[15: 8], o21_22[111:104], o21_22[79:72], o21_22[47:40], o21_22[15: 8], o21_23[111:104], o21_23[79:72], o21_23[47:40], o21_23[15: 8] };
		i33_03 <= { o22_20[103: 96], o22_20[71:64], o22_20[39:32], o22_20[ 7: 0], o22_21[103: 96], o22_21[71:64], o22_21[39:32], o22_21[ 7: 0], o22_22[103: 96], o22_22[71:64], o22_22[39:32], o22_22[ 7: 0], o22_23[103: 96], o22_23[71:64], o22_23[39:32], o22_23[ 7: 0] }; 

		i33_10 <= { o33_00[127:108], o33_00[107:96] ^ 12'h023C, o33_00[95:0] };
		i33_11 <= { o33_01[127:108], o33_01[107:96] ^ 12'h0231, o33_01[95:0] };
		i33_12 <= { o33_02[127:108], o33_02[107:96] ^ 12'h0236, o33_02[95:0] };
		i33_13 <= { o33_03[127:108], o33_03[107:96] ^ 12'h023B, o33_03[95:0] };

		i33_20 <= { o33_10[127:120], o33_11[127:120], o33_12[127:120], o33_13[127:120], o33_10[119:112], o33_11[119:112], o33_12[119:112], o33_13[119:112], o33_10[111:104], o33_11[111:104], o33_12[111:104], o33_13[111:104], o33_10[103: 96], o33_11[103: 96], o33_12[103: 96], o33_13[103: 96] };
		i33_21 <= { o33_10[ 95: 88], o33_11[ 95: 88], o33_12[ 95: 88], o33_13[ 95: 88], o33_10[ 87: 80], o33_11[ 87: 80], o33_12[ 87: 80], o33_13[ 87: 80], o33_10[ 79: 72], o33_11[ 79: 72], o33_12[ 79: 72], o33_13[ 79: 72],	o33_10[ 71: 64], o33_11[ 71: 64], o33_12[ 71: 64], o33_13[ 71: 64] };
		i33_22 <= { o33_10[ 63: 56], o33_11[ 63: 56], o33_12[ 63: 56], o33_13[ 63: 56], o33_10[ 55: 48], o33_11[ 55: 48], o33_12[ 55: 48], o33_13[ 55: 48], o33_10[ 47: 40], o33_11[ 47: 40], o33_12[ 47: 40], o33_13[ 47: 40], o33_10[ 39: 32], o33_11[ 39: 32], o33_12[ 39: 32], o33_13[ 39: 32] };
		i33_23 <= { o33_10[ 31: 24], o33_11[ 31: 24], o33_12[ 31: 24], o33_13[ 31: 24], o33_10[ 23: 16], o33_11[ 23: 16], o33_12[ 23: 16], o33_13[ 23: 16], o33_10[ 15:  8], o33_11[ 15:  8], o33_12[ 15:  8], o33_13[ 15:  8], o33_10[  7:  0], o33_11[  7:  0], o33_12[  7:  0], o33_13[  7:  0] };

	end

	// ROUND 4

	reg  [127:0] i40_00, i40_01, i40_02, i40_03, i40_10, i40_11, i40_12, i40_13, i40_20, i40_21, i40_22, i40_23;
	wire [127:0] o40_00, o40_01, o40_02, o40_03, o40_10, o40_11, o40_12, o40_13, o40_20, o40_21, o40_22, o40_23;

	aes_round r40_00 (clk, i40_00, o40_00);
	aes_round r40_01 (clk, i40_01, o40_01);
	aes_round r40_02 (clk, i40_02, o40_02);
	aes_round r40_03 (clk, i40_03, o40_03);

	aes_round r40_10 (clk, i40_10, o40_10);
	aes_round r40_11 (clk, i40_11, o40_11);
	aes_round r40_12 (clk, i40_12, o40_12);
	aes_round r40_13 (clk, i40_13, o40_13);
	
	echo_mix  r40_20 (clk, i40_20, o40_20);
	echo_mix  r40_21 (clk, i40_21, o40_21);
	echo_mix  r40_22 (clk, i40_22, o40_22);
	echo_mix  r40_23 (clk, i40_23, o40_23);

	always @ ( posedge clk ) begin

		i40_00 <= { o30_20[127:120], o30_20[95:88], o30_20[63:56], o30_20[31:24], o30_21[127:120], o30_21[95:88], o30_21[63:56], o30_21[31:24], o30_22[127:120], o30_22[95:88], o30_22[63:56], o30_22[31:24], o30_23[127:120], o30_23[95:88], o30_23[63:56], o30_23[31:24] };
		i40_01 <= { o31_20[119:112], o31_20[87:80], o31_20[55:48], o31_20[23:16], o31_21[119:112], o31_21[87:80], o31_21[55:48], o31_21[23:16], o31_22[119:112], o31_22[87:80], o31_22[55:48], o31_22[23:16], o31_23[119:112], o31_23[87:80], o31_23[55:48], o31_23[23:16] };
		i40_02 <= { o32_20[111:104], o32_20[79:72], o32_20[47:40], o32_20[15: 8], o32_21[111:104], o32_21[79:72], o32_21[47:40], o32_21[15: 8], o32_22[111:104], o32_22[79:72], o32_22[47:40], o32_22[15: 8], o32_23[111:104], o32_23[79:72], o32_23[47:40], o32_23[15: 8] };
		i40_03 <= { o33_20[103: 96], o33_20[71:64], o33_20[39:32], o33_20[ 7: 0], o33_21[103: 96], o33_21[71:64], o33_21[39:32], o33_21[ 7: 0], o33_22[103: 96], o33_22[71:64], o33_22[39:32], o33_22[ 7: 0], o33_23[103: 96], o33_23[71:64], o33_23[39:32], o33_23[ 7: 0] }; 

		i40_10 <= { o40_00[127:108], o40_00[107:96] ^ 12'h0240, o40_00[95:0] };
		i40_11 <= { o40_01[127:108], o40_01[107:96] ^ 12'h0245, o40_01[95:0] };
		i40_12 <= { o40_02[127:108], o40_02[107:96] ^ 12'h024A, o40_02[95:0] };
		i40_13 <= { o40_03[127:108], o40_03[107:96] ^ 12'h024F, o40_03[95:0] };

		i40_20 <= { o40_10[127:120], o40_11[127:120], o40_12[127:120], o40_13[127:120], o40_10[119:112], o40_11[119:112], o40_12[119:112], o40_13[119:112], o40_10[111:104], o40_11[111:104], o40_12[111:104], o40_13[111:104], o40_10[103: 96], o40_11[103: 96], o40_12[103: 96], o40_13[103: 96] };
		i40_21 <= { o40_10[ 95: 88], o40_11[ 95: 88], o40_12[ 95: 88], o40_13[ 95: 88], o40_10[ 87: 80], o40_11[ 87: 80], o40_12[ 87: 80], o40_13[ 87: 80], o40_10[ 79: 72], o40_11[ 79: 72], o40_12[ 79: 72], o40_13[ 79: 72],	o40_10[ 71: 64], o40_11[ 71: 64], o40_12[ 71: 64], o40_13[ 71: 64] };
		i40_22 <= { o40_10[ 63: 56], o40_11[ 63: 56], o40_12[ 63: 56], o40_13[ 63: 56], o40_10[ 55: 48], o40_11[ 55: 48], o40_12[ 55: 48], o40_13[ 55: 48], o40_10[ 47: 40], o40_11[ 47: 40], o40_12[ 47: 40], o40_13[ 47: 40], o40_10[ 39: 32], o40_11[ 39: 32], o40_12[ 39: 32], o40_13[ 39: 32] };
		i40_23 <= { o40_10[ 31: 24], o40_11[ 31: 24], o40_12[ 31: 24], o40_13[ 31: 24], o40_10[ 23: 16], o40_11[ 23: 16], o40_12[ 23: 16], o40_13[ 23: 16], o40_10[ 15:  8], o40_11[ 15:  8], o40_12[ 15:  8], o40_13[ 15:  8], o40_10[  7:  0], o40_11[  7:  0], o40_12[  7:  0], o40_13[  7:  0] };
		
	end

	reg  [127:0] i41_00, i41_01, i41_02, i41_03, i41_10, i41_11, i41_12, i41_13, i41_20, i41_21, i41_22, i41_23;
	wire [127:0] o41_00, o41_01, o41_02, o41_03, o41_10, o41_11, o41_12, o41_13, o41_20, o41_21, o41_22, o41_23;

	aes_round r41_00 (clk, i41_00, o41_00);
	aes_round r41_01 (clk, i41_01, o41_01);
	aes_round r41_02 (clk, i41_02, o41_02);
	aes_round r41_03 (clk, i41_03, o41_03);

	aes_round r41_10 (clk, i41_10, o41_10);
	aes_round r41_11 (clk, i41_11, o41_11);
	aes_round r41_12 (clk, i41_12, o41_12);
	aes_round r41_13 (clk, i41_13, o41_13);
	
	echo_mix  r41_20 (clk, i41_20, o41_20);
	echo_mix  r41_21 (clk, i41_21, o41_21);
	echo_mix  r41_22 (clk, i41_22, o41_22);
	echo_mix  r41_23 (clk, i41_23, o41_23);

	always @ ( posedge clk ) begin

		i41_00 <= { o31_20[127:120], o31_20[95:88], o31_20[63:56], o31_20[31:24], o31_21[127:120], o31_21[95:88], o31_21[63:56], o31_21[31:24], o31_22[127:120], o31_22[95:88], o31_22[63:56], o31_22[31:24], o31_23[127:120], o31_23[95:88], o31_23[63:56], o31_23[31:24] };
		i41_01 <= { o32_20[119:112], o32_20[87:80], o32_20[55:48], o32_20[23:16], o32_21[119:112], o32_21[87:80], o32_21[55:48], o32_21[23:16], o32_22[119:112], o32_22[87:80], o32_22[55:48], o32_22[23:16], o32_23[119:112], o32_23[87:80], o32_23[55:48], o32_23[23:16] };
		i41_02 <= { o33_20[111:104], o33_20[79:72], o33_20[47:40], o33_20[15: 8], o33_21[111:104], o33_21[79:72], o33_21[47:40], o33_21[15: 8], o33_22[111:104], o33_22[79:72], o33_22[47:40], o33_22[15: 8], o33_23[111:104], o33_23[79:72], o33_23[47:40], o33_23[15: 8] };
		i41_03 <= { o30_20[103: 96], o30_20[71:64], o30_20[39:32], o30_20[ 7: 0], o30_21[103: 96], o30_21[71:64], o30_21[39:32], o30_21[ 7: 0], o30_22[103: 96], o30_22[71:64], o30_22[39:32], o30_22[ 7: 0], o30_23[103: 96], o30_23[71:64], o30_23[39:32], o30_23[ 7: 0] };

		i41_10 <= { o41_00[127:108], o41_00[107:96] ^ 12'h0244, o41_00[95:0] };
		i41_11 <= { o41_01[127:108], o41_01[107:96] ^ 12'h0249, o41_01[95:0] };
		i41_12 <= { o41_02[127:108], o41_02[107:96] ^ 12'h024E, o41_02[95:0] };
		i41_13 <= { o41_03[127:108], o41_03[107:96] ^ 12'h0243, o41_03[95:0] };

		i41_20 <= { o41_10[127:120], o41_11[127:120], o41_12[127:120], o41_13[127:120], o41_10[119:112], o41_11[119:112], o41_12[119:112], o41_13[119:112], o41_10[111:104], o41_11[111:104], o41_12[111:104], o41_13[111:104], o41_10[103: 96], o41_11[103: 96], o41_12[103: 96], o41_13[103: 96] };
		i41_21 <= { o41_10[ 95: 88], o41_11[ 95: 88], o41_12[ 95: 88], o41_13[ 95: 88], o41_10[ 87: 80], o41_11[ 87: 80], o41_12[ 87: 80], o41_13[ 87: 80], o41_10[ 79: 72], o41_11[ 79: 72], o41_12[ 79: 72], o41_13[ 79: 72],	o41_10[ 71: 64], o41_11[ 71: 64], o41_12[ 71: 64], o41_13[ 71: 64] };
		i41_22 <= { o41_10[ 63: 56], o41_11[ 63: 56], o41_12[ 63: 56], o41_13[ 63: 56], o41_10[ 55: 48], o41_11[ 55: 48], o41_12[ 55: 48], o41_13[ 55: 48], o41_10[ 47: 40], o41_11[ 47: 40], o41_12[ 47: 40], o41_13[ 47: 40], o41_10[ 39: 32], o41_11[ 39: 32], o41_12[ 39: 32], o41_13[ 39: 32] };
		i41_23 <= { o41_10[ 31: 24], o41_11[ 31: 24], o41_12[ 31: 24], o41_13[ 31: 24], o41_10[ 23: 16], o41_11[ 23: 16], o41_12[ 23: 16], o41_13[ 23: 16], o41_10[ 15:  8], o41_11[ 15:  8], o41_12[ 15:  8], o41_13[ 15:  8], o41_10[  7:  0], o41_11[  7:  0], o41_12[  7:  0], o41_13[  7:  0] };

	end

	reg  [127:0] i42_00, i42_01, i42_02, i42_03, i42_10, i42_11, i42_12, i42_13, i42_20, i42_21, i42_22, i42_23;
	wire [127:0] o42_00, o42_01, o42_02, o42_03, o42_10, o42_11, o42_12, o42_13, o42_20, o42_21, o42_22, o42_23;

	aes_round r42_00 (clk, i42_00, o42_00);
	aes_round r42_01 (clk, i42_01, o42_01);
	aes_round r42_02 (clk, i42_02, o42_02);
	aes_round r42_03 (clk, i42_03, o42_03);

	aes_round r42_10 (clk, i42_10, o42_10);
	aes_round r42_11 (clk, i42_11, o42_11);
	aes_round r42_12 (clk, i42_12, o42_12);
	aes_round r42_13 (clk, i42_13, o42_13);
	
	echo_mix  r42_20 (clk, i42_20, o42_20);
	echo_mix  r42_21 (clk, i42_21, o42_21);
	echo_mix  r42_22 (clk, i42_22, o42_22);
	echo_mix  r42_23 (clk, i42_23, o42_23);

	always @ ( posedge clk ) begin

		i42_00 <= { o32_20[127:120], o32_20[95:88], o32_20[63:56], o32_20[31:24], o32_21[127:120], o32_21[95:88], o32_21[63:56], o32_21[31:24], o32_22[127:120], o32_22[95:88], o32_22[63:56], o32_22[31:24], o32_23[127:120], o32_23[95:88], o32_23[63:56], o32_23[31:24] };
		i42_01 <= { o33_20[119:112], o33_20[87:80], o33_20[55:48], o33_20[23:16], o33_21[119:112], o33_21[87:80], o33_21[55:48], o33_21[23:16], o33_22[119:112], o33_22[87:80], o33_22[55:48], o33_22[23:16], o33_23[119:112], o33_23[87:80], o33_23[55:48], o33_23[23:16] };
		i42_02 <= { o30_20[111:104], o30_20[79:72], o30_20[47:40], o30_20[15: 8], o30_21[111:104], o30_21[79:72], o30_21[47:40], o30_21[15: 8], o30_22[111:104], o30_22[79:72], o30_22[47:40], o30_22[15: 8], o30_23[111:104], o30_23[79:72], o30_23[47:40], o30_23[15: 8] };
		i42_03 <= { o31_20[103: 96], o31_20[71:64], o31_20[39:32], o31_20[ 7: 0], o31_21[103: 96], o31_21[71:64], o31_21[39:32], o31_21[ 7: 0], o31_22[103: 96], o31_22[71:64], o31_22[39:32], o31_22[ 7: 0], o31_23[103: 96], o31_23[71:64], o31_23[39:32], o31_23[ 7: 0] }; 

		i42_10 <= { o42_00[127:108], o42_00[107:96] ^ 12'h0248, o42_00[95:0] };
		i42_11 <= { o42_01[127:108], o42_01[107:96] ^ 12'h024D, o42_01[95:0] };
		i42_12 <= { o42_02[127:108], o42_02[107:96] ^ 12'h0242, o42_02[95:0] };
		i42_13 <= { o42_03[127:108], o42_03[107:96] ^ 12'h0247, o42_03[95:0] };

		i42_20 <= { o42_10[127:120], o42_11[127:120], o42_12[127:120], o42_13[127:120], o42_10[119:112], o42_11[119:112], o42_12[119:112], o42_13[119:112], o42_10[111:104], o42_11[111:104], o42_12[111:104], o42_13[111:104], o42_10[103: 96], o42_11[103: 96], o42_12[103: 96], o42_13[103: 96] };
		i42_21 <= { o42_10[ 95: 88], o42_11[ 95: 88], o42_12[ 95: 88], o42_13[ 95: 88], o42_10[ 87: 80], o42_11[ 87: 80], o42_12[ 87: 80], o42_13[ 87: 80], o42_10[ 79: 72], o42_11[ 79: 72], o42_12[ 79: 72], o42_13[ 79: 72],	o42_10[ 71: 64], o42_11[ 71: 64], o42_12[ 71: 64], o42_13[ 71: 64] };
		i42_22 <= { o42_10[ 63: 56], o42_11[ 63: 56], o42_12[ 63: 56], o42_13[ 63: 56], o42_10[ 55: 48], o42_11[ 55: 48], o42_12[ 55: 48], o42_13[ 55: 48], o42_10[ 47: 40], o42_11[ 47: 40], o42_12[ 47: 40], o42_13[ 47: 40], o42_10[ 39: 32], o42_11[ 39: 32], o42_12[ 39: 32], o42_13[ 39: 32] };
		i42_23 <= { o42_10[ 31: 24], o42_11[ 31: 24], o42_12[ 31: 24], o42_13[ 31: 24], o42_10[ 23: 16], o42_11[ 23: 16], o42_12[ 23: 16], o42_13[ 23: 16], o42_10[ 15:  8], o42_11[ 15:  8], o42_12[ 15:  8], o42_13[ 15:  8], o42_10[  7:  0], o42_11[  7:  0], o42_12[  7:  0], o42_13[  7:  0] };

	end

	reg  [127:0] i43_00, i43_01, i43_02, i43_03, i43_10, i43_11, i43_12, i43_13, i43_20, i43_21, i43_22, i43_23;
	wire [127:0] o43_00, o43_01, o43_02, o43_03, o43_10, o43_11, o43_12, o43_13, o43_20, o43_21, o43_22, o43_23;

	aes_round r43_00 (clk, i43_00, o43_00);
	aes_round r43_01 (clk, i43_01, o43_01);
	aes_round r43_02 (clk, i43_02, o43_02);
	aes_round r43_03 (clk, i43_03, o43_03);

	aes_round r43_10 (clk, i43_10, o43_10);
	aes_round r43_11 (clk, i43_11, o43_11);
	aes_round r43_12 (clk, i43_12, o43_12);
	aes_round r43_13 (clk, i43_13, o43_13);
	
	echo_mix  r43_20 (clk, i43_20, o43_20);
	echo_mix  r43_21 (clk, i43_21, o43_21);
	echo_mix  r43_22 (clk, i43_22, o43_22);
	echo_mix  r43_23 (clk, i43_23, o43_23);

	always @ ( posedge clk ) begin

		i43_00 <= { o33_20[127:120], o33_20[95:88], o33_20[63:56], o33_20[31:24], o33_21[127:120], o33_21[95:88], o33_21[63:56], o33_21[31:24], o33_22[127:120], o33_22[95:88], o33_22[63:56], o33_22[31:24], o33_23[127:120], o33_23[95:88], o33_23[63:56], o33_23[31:24] };
		i43_01 <= { o30_20[119:112], o30_20[87:80], o30_20[55:48], o30_20[23:16], o30_21[119:112], o30_21[87:80], o30_21[55:48], o30_21[23:16], o30_22[119:112], o30_22[87:80], o30_22[55:48], o30_22[23:16], o30_23[119:112], o30_23[87:80], o30_23[55:48], o30_23[23:16] };
		i43_02 <= { o31_20[111:104], o31_20[79:72], o31_20[47:40], o31_20[15: 8], o31_21[111:104], o31_21[79:72], o31_21[47:40], o31_21[15: 8], o31_22[111:104], o31_22[79:72], o31_22[47:40], o31_22[15: 8], o31_23[111:104], o31_23[79:72], o31_23[47:40], o31_23[15: 8] };
		i43_03 <= { o32_20[103: 96], o32_20[71:64], o32_20[39:32], o32_20[ 7: 0], o32_21[103: 96], o32_21[71:64], o32_21[39:32], o32_21[ 7: 0], o32_22[103: 96], o32_22[71:64], o32_22[39:32], o32_22[ 7: 0], o32_23[103: 96], o32_23[71:64], o32_23[39:32], o32_23[ 7: 0] }; 

		i43_10 <= { o43_00[127:108], o43_00[107:96] ^ 12'h024C, o43_00[95:0] };
		i43_11 <= { o43_01[127:108], o43_01[107:96] ^ 12'h0241, o43_01[95:0] };
		i43_12 <= { o43_02[127:108], o43_02[107:96] ^ 12'h0246, o43_02[95:0] };
		i43_13 <= { o43_03[127:108], o43_03[107:96] ^ 12'h024B, o43_03[95:0] };

		i43_20 <= { o43_10[127:120], o43_11[127:120], o43_12[127:120], o43_13[127:120], o43_10[119:112], o43_11[119:112], o43_12[119:112], o43_13[119:112], o43_10[111:104], o43_11[111:104], o43_12[111:104], o43_13[111:104], o43_10[103: 96], o43_11[103: 96], o43_12[103: 96], o43_13[103: 96] };
		i43_21 <= { o43_10[ 95: 88], o43_11[ 95: 88], o43_12[ 95: 88], o43_13[ 95: 88], o43_10[ 87: 80], o43_11[ 87: 80], o43_12[ 87: 80], o43_13[ 87: 80], o43_10[ 79: 72], o43_11[ 79: 72], o43_12[ 79: 72], o43_13[ 79: 72],	o43_10[ 71: 64], o43_11[ 71: 64], o43_12[ 71: 64], o43_13[ 71: 64] };
		i43_22 <= { o43_10[ 63: 56], o43_11[ 63: 56], o43_12[ 63: 56], o43_13[ 63: 56], o43_10[ 55: 48], o43_11[ 55: 48], o43_12[ 55: 48], o43_13[ 55: 48], o43_10[ 47: 40], o43_11[ 47: 40], o43_12[ 47: 40], o43_13[ 47: 40], o43_10[ 39: 32], o43_11[ 39: 32], o43_12[ 39: 32], o43_13[ 39: 32] };
		i43_23 <= { o43_10[ 31: 24], o43_11[ 31: 24], o43_12[ 31: 24], o43_13[ 31: 24], o43_10[ 23: 16], o43_11[ 23: 16], o43_12[ 23: 16], o43_13[ 23: 16], o43_10[ 15:  8], o43_11[ 15:  8], o43_12[ 15:  8], o43_13[ 15:  8], o43_10[  7:  0], o43_11[  7:  0], o43_12[  7:  0], o43_13[  7:  0] };

	end

	// ROUND 5

	reg  [127:0] i50_00, i50_01, i50_02, i50_03, i50_10, i50_11, i50_12, i50_13, i50_20, i50_21, i50_22, i50_23;
	wire [127:0] o50_00, o50_01, o50_02, o50_03, o50_10, o50_11, o50_12, o50_13, o50_20, o50_21, o50_22, o50_23;

	aes_round r50_00 (clk, i50_00, o50_00);
	aes_round r50_01 (clk, i50_01, o50_01);
	aes_round r50_02 (clk, i50_02, o50_02);
	aes_round r50_03 (clk, i50_03, o50_03);

	aes_round r50_10 (clk, i50_10, o50_10);
	aes_round r50_11 (clk, i50_11, o50_11);
	aes_round r50_12 (clk, i50_12, o50_12);
	aes_round r50_13 (clk, i50_13, o50_13);
	
	echo_mix  r50_20 (clk, i50_20, o50_20);
	echo_mix  r50_21 (clk, i50_21, o50_21);
	echo_mix  r50_22 (clk, i50_22, o50_22);
	echo_mix  r50_23 (clk, i50_23, o50_23);

	always @ ( posedge clk ) begin

		i50_00 <= { o40_20[127:120], o40_20[95:88], o40_20[63:56], o40_20[31:24], o40_21[127:120], o40_21[95:88], o40_21[63:56], o40_21[31:24], o40_22[127:120], o40_22[95:88], o40_22[63:56], o40_22[31:24], o40_23[127:120], o40_23[95:88], o40_23[63:56], o40_23[31:24] };
		i50_01 <= { o41_20[119:112], o41_20[87:80], o41_20[55:48], o41_20[23:16], o41_21[119:112], o41_21[87:80], o41_21[55:48], o41_21[23:16], o41_22[119:112], o41_22[87:80], o41_22[55:48], o41_22[23:16], o41_23[119:112], o41_23[87:80], o41_23[55:48], o41_23[23:16] };
		i50_02 <= { o42_20[111:104], o42_20[79:72], o42_20[47:40], o42_20[15: 8], o42_21[111:104], o42_21[79:72], o42_21[47:40], o42_21[15: 8], o42_22[111:104], o42_22[79:72], o42_22[47:40], o42_22[15: 8], o42_23[111:104], o42_23[79:72], o42_23[47:40], o42_23[15: 8] };
		i50_03 <= { o43_20[103: 96], o43_20[71:64], o43_20[39:32], o43_20[ 7: 0], o43_21[103: 96], o43_21[71:64], o43_21[39:32], o43_21[ 7: 0], o43_22[103: 96], o43_22[71:64], o43_22[39:32], o43_22[ 7: 0], o43_23[103: 96], o43_23[71:64], o43_23[39:32], o43_23[ 7: 0] }; 

		i50_10 <= { o50_00[127:108], o50_00[107:96] ^ 12'h0250, o50_00[95:0] };
		i50_11 <= { o50_01[127:108], o50_01[107:96] ^ 12'h0255, o50_01[95:0] };
		i50_12 <= { o50_02[127:108], o50_02[107:96] ^ 12'h025A, o50_02[95:0] };
		i50_13 <= { o50_03[127:108], o50_03[107:96] ^ 12'h025F, o50_03[95:0] };

		i50_20 <= { o50_10[127:120], o50_11[127:120], o50_12[127:120], o50_13[127:120], o50_10[119:112], o50_11[119:112], o50_12[119:112], o50_13[119:112], o50_10[111:104], o50_11[111:104], o50_12[111:104], o50_13[111:104], o50_10[103: 96], o50_11[103: 96], o50_12[103: 96], o50_13[103: 96] };
		i50_21 <= { o50_10[ 95: 88], o50_11[ 95: 88], o50_12[ 95: 88], o50_13[ 95: 88], o50_10[ 87: 80], o50_11[ 87: 80], o50_12[ 87: 80], o50_13[ 87: 80], o50_10[ 79: 72], o50_11[ 79: 72], o50_12[ 79: 72], o50_13[ 79: 72],	o50_10[ 71: 64], o50_11[ 71: 64], o50_12[ 71: 64], o50_13[ 71: 64] };
		i50_22 <= { o50_10[ 63: 56], o50_11[ 63: 56], o50_12[ 63: 56], o50_13[ 63: 56], o50_10[ 55: 48], o50_11[ 55: 48], o50_12[ 55: 48], o50_13[ 55: 48], o50_10[ 47: 40], o50_11[ 47: 40], o50_12[ 47: 40], o50_13[ 47: 40], o50_10[ 39: 32], o50_11[ 39: 32], o50_12[ 39: 32], o50_13[ 39: 32] };
		i50_23 <= { o50_10[ 31: 24], o50_11[ 31: 24], o50_12[ 31: 24], o50_13[ 31: 24], o50_10[ 23: 16], o50_11[ 23: 16], o50_12[ 23: 16], o50_13[ 23: 16], o50_10[ 15:  8], o50_11[ 15:  8], o50_12[ 15:  8], o50_13[ 15:  8], o50_10[  7:  0], o50_11[  7:  0], o50_12[  7:  0], o50_13[  7:  0] };
		
	end

	reg  [127:0] i51_00, i51_01, i51_02, i51_03, i51_10, i51_11, i51_12, i51_13, i51_20, i51_21, i51_22, i51_23;
	wire [127:0] o51_00, o51_01, o51_02, o51_03, o51_10, o51_11, o51_12, o51_13, o51_20, o51_21, o51_22, o51_23;

	aes_round r51_00 (clk, i51_00, o51_00);
	aes_round r51_01 (clk, i51_01, o51_01);
	aes_round r51_02 (clk, i51_02, o51_02);
	aes_round r51_03 (clk, i51_03, o51_03);

	aes_round r51_10 (clk, i51_10, o51_10);
	aes_round r51_11 (clk, i51_11, o51_11);
	aes_round r51_12 (clk, i51_12, o51_12);
	aes_round r51_13 (clk, i51_13, o51_13);
	
	echo_mix  r51_20 (clk, i51_20, o51_20);
	echo_mix  r51_21 (clk, i51_21, o51_21);
	echo_mix  r51_22 (clk, i51_22, o51_22);
	echo_mix  r51_23 (clk, i51_23, o51_23);

	always @ ( posedge clk ) begin

		i51_00 <= { o41_20[127:120], o41_20[95:88], o41_20[63:56], o41_20[31:24], o41_21[127:120], o41_21[95:88], o41_21[63:56], o41_21[31:24], o41_22[127:120], o41_22[95:88], o41_22[63:56], o41_22[31:24], o41_23[127:120], o41_23[95:88], o41_23[63:56], o41_23[31:24] };
		i51_01 <= { o42_20[119:112], o42_20[87:80], o42_20[55:48], o42_20[23:16], o42_21[119:112], o42_21[87:80], o42_21[55:48], o42_21[23:16], o42_22[119:112], o42_22[87:80], o42_22[55:48], o42_22[23:16], o42_23[119:112], o42_23[87:80], o42_23[55:48], o42_23[23:16] };
		i51_02 <= { o43_20[111:104], o43_20[79:72], o43_20[47:40], o43_20[15: 8], o43_21[111:104], o43_21[79:72], o43_21[47:40], o43_21[15: 8], o43_22[111:104], o43_22[79:72], o43_22[47:40], o43_22[15: 8], o43_23[111:104], o43_23[79:72], o43_23[47:40], o43_23[15: 8] };
		i51_03 <= { o40_20[103: 96], o40_20[71:64], o40_20[39:32], o40_20[ 7: 0], o40_21[103: 96], o40_21[71:64], o40_21[39:32], o40_21[ 7: 0], o40_22[103: 96], o40_22[71:64], o40_22[39:32], o40_22[ 7: 0], o40_23[103: 96], o40_23[71:64], o40_23[39:32], o40_23[ 7: 0] };

		i51_10 <= { o51_00[127:108], o51_00[107:96] ^ 12'h0254, o51_00[95:0] };
		i51_11 <= { o51_01[127:108], o51_01[107:96] ^ 12'h0259, o51_01[95:0] };
		i51_12 <= { o51_02[127:108], o51_02[107:96] ^ 12'h025E, o51_02[95:0] };
		i51_13 <= { o51_03[127:108], o51_03[107:96] ^ 12'h0253, o51_03[95:0] };

		i51_20 <= { o51_10[127:120], o51_11[127:120], o51_12[127:120], o51_13[127:120], o51_10[119:112], o51_11[119:112], o51_12[119:112], o51_13[119:112], o51_10[111:104], o51_11[111:104], o51_12[111:104], o51_13[111:104], o51_10[103: 96], o51_11[103: 96], o51_12[103: 96], o51_13[103: 96] };
		i51_21 <= { o51_10[ 95: 88], o51_11[ 95: 88], o51_12[ 95: 88], o51_13[ 95: 88], o51_10[ 87: 80], o51_11[ 87: 80], o51_12[ 87: 80], o51_13[ 87: 80], o51_10[ 79: 72], o51_11[ 79: 72], o51_12[ 79: 72], o51_13[ 79: 72],	o51_10[ 71: 64], o51_11[ 71: 64], o51_12[ 71: 64], o51_13[ 71: 64] };
		i51_22 <= { o51_10[ 63: 56], o51_11[ 63: 56], o51_12[ 63: 56], o51_13[ 63: 56], o51_10[ 55: 48], o51_11[ 55: 48], o51_12[ 55: 48], o51_13[ 55: 48], o51_10[ 47: 40], o51_11[ 47: 40], o51_12[ 47: 40], o51_13[ 47: 40], o51_10[ 39: 32], o51_11[ 39: 32], o51_12[ 39: 32], o51_13[ 39: 32] };
		i51_23 <= { o51_10[ 31: 24], o51_11[ 31: 24], o51_12[ 31: 24], o51_13[ 31: 24], o51_10[ 23: 16], o51_11[ 23: 16], o51_12[ 23: 16], o51_13[ 23: 16], o51_10[ 15:  8], o51_11[ 15:  8], o51_12[ 15:  8], o51_13[ 15:  8], o51_10[  7:  0], o51_11[  7:  0], o51_12[  7:  0], o51_13[  7:  0] };

	end

	reg  [127:0] i52_00, i52_01, i52_02, i52_03, i52_10, i52_11, i52_12, i52_13, i52_20, i52_21, i52_22, i52_23;
	wire [127:0] o52_00, o52_01, o52_02, o52_03, o52_10, o52_11, o52_12, o52_13, o52_20, o52_21, o52_22, o52_23;

	aes_round r52_00 (clk, i52_00, o52_00);
	aes_round r52_01 (clk, i52_01, o52_01);
	aes_round r52_02 (clk, i52_02, o52_02);
	aes_round r52_03 (clk, i52_03, o52_03);

	aes_round r52_10 (clk, i52_10, o52_10);
	aes_round r52_11 (clk, i52_11, o52_11);
	aes_round r52_12 (clk, i52_12, o52_12);
	aes_round r52_13 (clk, i52_13, o52_13);
	
	echo_mix  r52_20 (clk, i52_20, o52_20);
	echo_mix  r52_21 (clk, i52_21, o52_21);
	echo_mix  r52_22 (clk, i52_22, o52_22);
	echo_mix  r52_23 (clk, i52_23, o52_23);

	always @ ( posedge clk ) begin

		i52_00 <= { o42_20[127:120], o42_20[95:88], o42_20[63:56], o42_20[31:24], o42_21[127:120], o42_21[95:88], o42_21[63:56], o42_21[31:24], o42_22[127:120], o42_22[95:88], o42_22[63:56], o42_22[31:24], o42_23[127:120], o42_23[95:88], o42_23[63:56], o42_23[31:24] };
		i52_01 <= { o43_20[119:112], o43_20[87:80], o43_20[55:48], o43_20[23:16], o43_21[119:112], o43_21[87:80], o43_21[55:48], o43_21[23:16], o43_22[119:112], o43_22[87:80], o43_22[55:48], o43_22[23:16], o43_23[119:112], o43_23[87:80], o43_23[55:48], o43_23[23:16] };
		i52_02 <= { o40_20[111:104], o40_20[79:72], o40_20[47:40], o40_20[15: 8], o40_21[111:104], o40_21[79:72], o40_21[47:40], o40_21[15: 8], o40_22[111:104], o40_22[79:72], o40_22[47:40], o40_22[15: 8], o40_23[111:104], o40_23[79:72], o40_23[47:40], o40_23[15: 8] };
		i52_03 <= { o41_20[103: 96], o41_20[71:64], o41_20[39:32], o41_20[ 7: 0], o41_21[103: 96], o41_21[71:64], o41_21[39:32], o41_21[ 7: 0], o41_22[103: 96], o41_22[71:64], o41_22[39:32], o41_22[ 7: 0], o41_23[103: 96], o41_23[71:64], o41_23[39:32], o41_23[ 7: 0] }; 

		i52_10 <= { o52_00[127:108], o52_00[107:96] ^ 12'h0258, o52_00[95:0] };
		i52_11 <= { o52_01[127:108], o52_01[107:96] ^ 12'h025D, o52_01[95:0] };
		i52_12 <= { o52_02[127:108], o52_02[107:96] ^ 12'h0252, o52_02[95:0] };
		i52_13 <= { o52_03[127:108], o52_03[107:96] ^ 12'h0257, o52_03[95:0] };

		i52_20 <= { o52_10[127:120], o52_11[127:120], o52_12[127:120], o52_13[127:120], o52_10[119:112], o52_11[119:112], o52_12[119:112], o52_13[119:112], o52_10[111:104], o52_11[111:104], o52_12[111:104], o52_13[111:104], o52_10[103: 96], o52_11[103: 96], o52_12[103: 96], o52_13[103: 96] };
		i52_21 <= { o52_10[ 95: 88], o52_11[ 95: 88], o52_12[ 95: 88], o52_13[ 95: 88], o52_10[ 87: 80], o52_11[ 87: 80], o52_12[ 87: 80], o52_13[ 87: 80], o52_10[ 79: 72], o52_11[ 79: 72], o52_12[ 79: 72], o52_13[ 79: 72],	o52_10[ 71: 64], o52_11[ 71: 64], o52_12[ 71: 64], o52_13[ 71: 64] };
		i52_22 <= { o52_10[ 63: 56], o52_11[ 63: 56], o52_12[ 63: 56], o52_13[ 63: 56], o52_10[ 55: 48], o52_11[ 55: 48], o52_12[ 55: 48], o52_13[ 55: 48], o52_10[ 47: 40], o52_11[ 47: 40], o52_12[ 47: 40], o52_13[ 47: 40], o52_10[ 39: 32], o52_11[ 39: 32], o52_12[ 39: 32], o52_13[ 39: 32] };
		i52_23 <= { o52_10[ 31: 24], o52_11[ 31: 24], o52_12[ 31: 24], o52_13[ 31: 24], o52_10[ 23: 16], o52_11[ 23: 16], o52_12[ 23: 16], o52_13[ 23: 16], o52_10[ 15:  8], o52_11[ 15:  8], o52_12[ 15:  8], o52_13[ 15:  8], o52_10[  7:  0], o52_11[  7:  0], o52_12[  7:  0], o52_13[  7:  0] };

	end

	reg  [127:0] i53_00, i53_01, i53_02, i53_03, i53_10, i53_11, i53_12, i53_13, i53_20, i53_21, i53_22, i53_23;
	wire [127:0] o53_00, o53_01, o53_02, o53_03, o53_10, o53_11, o53_12, o53_13, o53_20, o53_21, o53_22, o53_23;

	aes_round r53_00 (clk, i53_00, o53_00);
	aes_round r53_01 (clk, i53_01, o53_01);
	aes_round r53_02 (clk, i53_02, o53_02);
	aes_round r53_03 (clk, i53_03, o53_03);

	aes_round r53_10 (clk, i53_10, o53_10);
	aes_round r53_11 (clk, i53_11, o53_11);
	aes_round r53_12 (clk, i53_12, o53_12);
	aes_round r53_13 (clk, i53_13, o53_13);
	
	echo_mix  r53_20 (clk, i53_20, o53_20);
	echo_mix  r53_21 (clk, i53_21, o53_21);
	echo_mix  r53_22 (clk, i53_22, o53_22);
	echo_mix  r53_23 (clk, i53_23, o53_23);

	always @ ( posedge clk ) begin

		i53_00 <= { o43_20[127:120], o43_20[95:88], o43_20[63:56], o43_20[31:24], o43_21[127:120], o43_21[95:88], o43_21[63:56], o43_21[31:24], o43_22[127:120], o43_22[95:88], o43_22[63:56], o43_22[31:24], o43_23[127:120], o43_23[95:88], o43_23[63:56], o43_23[31:24] };
		i53_01 <= { o40_20[119:112], o40_20[87:80], o40_20[55:48], o40_20[23:16], o40_21[119:112], o40_21[87:80], o40_21[55:48], o40_21[23:16], o40_22[119:112], o40_22[87:80], o40_22[55:48], o40_22[23:16], o40_23[119:112], o40_23[87:80], o40_23[55:48], o40_23[23:16] };
		i53_02 <= { o41_20[111:104], o41_20[79:72], o41_20[47:40], o41_20[15: 8], o41_21[111:104], o41_21[79:72], o41_21[47:40], o41_21[15: 8], o41_22[111:104], o41_22[79:72], o41_22[47:40], o41_22[15: 8], o41_23[111:104], o41_23[79:72], o41_23[47:40], o41_23[15: 8] };
		i53_03 <= { o42_20[103: 96], o42_20[71:64], o42_20[39:32], o42_20[ 7: 0], o42_21[103: 96], o42_21[71:64], o42_21[39:32], o42_21[ 7: 0], o42_22[103: 96], o42_22[71:64], o42_22[39:32], o42_22[ 7: 0], o42_23[103: 96], o42_23[71:64], o42_23[39:32], o42_23[ 7: 0] }; 

		i53_10 <= { o53_00[127:108], o53_00[107:96] ^ 12'h025C, o53_00[95:0] };
		i53_11 <= { o53_01[127:108], o53_01[107:96] ^ 12'h0251, o53_01[95:0] };
		i53_12 <= { o53_02[127:108], o53_02[107:96] ^ 12'h0256, o53_02[95:0] };
		i53_13 <= { o53_03[127:108], o53_03[107:96] ^ 12'h025B, o53_03[95:0] };

		i53_20 <= { o53_10[127:120], o53_11[127:120], o53_12[127:120], o53_13[127:120], o53_10[119:112], o53_11[119:112], o53_12[119:112], o53_13[119:112], o53_10[111:104], o53_11[111:104], o53_12[111:104], o53_13[111:104], o53_10[103: 96], o53_11[103: 96], o53_12[103: 96], o53_13[103: 96] };
		i53_21 <= { o53_10[ 95: 88], o53_11[ 95: 88], o53_12[ 95: 88], o53_13[ 95: 88], o53_10[ 87: 80], o53_11[ 87: 80], o53_12[ 87: 80], o53_13[ 87: 80], o53_10[ 79: 72], o53_11[ 79: 72], o53_12[ 79: 72], o53_13[ 79: 72],	o53_10[ 71: 64], o53_11[ 71: 64], o53_12[ 71: 64], o53_13[ 71: 64] };
		i53_22 <= { o53_10[ 63: 56], o53_11[ 63: 56], o53_12[ 63: 56], o53_13[ 63: 56], o53_10[ 55: 48], o53_11[ 55: 48], o53_12[ 55: 48], o53_13[ 55: 48], o53_10[ 47: 40], o53_11[ 47: 40], o53_12[ 47: 40], o53_13[ 47: 40], o53_10[ 39: 32], o53_11[ 39: 32], o53_12[ 39: 32], o53_13[ 39: 32] };
		i53_23 <= { o53_10[ 31: 24], o53_11[ 31: 24], o53_12[ 31: 24], o53_13[ 31: 24], o53_10[ 23: 16], o53_11[ 23: 16], o53_12[ 23: 16], o53_13[ 23: 16], o53_10[ 15:  8], o53_11[ 15:  8], o53_12[ 15:  8], o53_13[ 15:  8], o53_10[  7:  0], o53_11[  7:  0], o53_12[  7:  0], o53_13[  7:  0] };

	end

	// ROUND 6

	reg  [127:0] i60_00, i60_01, i60_02, i60_03, i60_10, i60_11, i60_12, i60_13, i60_20, i60_21, i60_22, i60_23;
	wire [127:0] o60_00, o60_01, o60_02, o60_03, o60_10, o60_11, o60_12, o60_13, o60_20, o60_21, o60_22, o60_23;

	aes_round r60_00 (clk, i60_00, o60_00);
	aes_round r60_01 (clk, i60_01, o60_01);
	aes_round r60_02 (clk, i60_02, o60_02);
	aes_round r60_03 (clk, i60_03, o60_03);

	aes_round r60_10 (clk, i60_10, o60_10);
	aes_round r60_11 (clk, i60_11, o60_11);
	aes_round r60_12 (clk, i60_12, o60_12);
	aes_round r60_13 (clk, i60_13, o60_13);
	
	echo_mix  r60_20 (clk, i60_20, o60_20);
	echo_mix  r60_21 (clk, i60_21, o60_21);
	echo_mix  r60_22 (clk, i60_22, o60_22);
	echo_mix  r60_23 (clk, i60_23, o60_23);

	always @ ( posedge clk ) begin

		i60_00 <= { o50_20[127:120], o50_20[95:88], o50_20[63:56], o50_20[31:24], o50_21[127:120], o50_21[95:88], o50_21[63:56], o50_21[31:24], o50_22[127:120], o50_22[95:88], o50_22[63:56], o50_22[31:24], o50_23[127:120], o50_23[95:88], o50_23[63:56], o50_23[31:24] };
		i60_01 <= { o51_20[119:112], o51_20[87:80], o51_20[55:48], o51_20[23:16], o51_21[119:112], o51_21[87:80], o51_21[55:48], o51_21[23:16], o51_22[119:112], o51_22[87:80], o51_22[55:48], o51_22[23:16], o51_23[119:112], o51_23[87:80], o51_23[55:48], o51_23[23:16] };
		i60_02 <= { o52_20[111:104], o52_20[79:72], o52_20[47:40], o52_20[15: 8], o52_21[111:104], o52_21[79:72], o52_21[47:40], o52_21[15: 8], o52_22[111:104], o52_22[79:72], o52_22[47:40], o52_22[15: 8], o52_23[111:104], o52_23[79:72], o52_23[47:40], o52_23[15: 8] };
		i60_03 <= { o53_20[103: 96], o53_20[71:64], o53_20[39:32], o53_20[ 7: 0], o53_21[103: 96], o53_21[71:64], o53_21[39:32], o53_21[ 7: 0], o53_22[103: 96], o53_22[71:64], o53_22[39:32], o53_22[ 7: 0], o53_23[103: 96], o53_23[71:64], o53_23[39:32], o53_23[ 7: 0] }; 

		i60_10 <= { o60_00[127:108], o60_00[107:96] ^ 12'h0260, o60_00[95:0] };
		i60_11 <= { o60_01[127:108], o60_01[107:96] ^ 12'h0265, o60_01[95:0] };
		i60_12 <= { o60_02[127:108], o60_02[107:96] ^ 12'h026A, o60_02[95:0] };
		i60_13 <= { o60_03[127:108], o60_03[107:96] ^ 12'h026F, o60_03[95:0] };

		i60_20 <= { o60_10[127:120], o60_11[127:120], o60_12[127:120], o60_13[127:120], o60_10[119:112], o60_11[119:112], o60_12[119:112], o60_13[119:112], o60_10[111:104], o60_11[111:104], o60_12[111:104], o60_13[111:104], o60_10[103: 96], o60_11[103: 96], o60_12[103: 96], o60_13[103: 96] };
		i60_21 <= { o60_10[ 95: 88], o60_11[ 95: 88], o60_12[ 95: 88], o60_13[ 95: 88], o60_10[ 87: 80], o60_11[ 87: 80], o60_12[ 87: 80], o60_13[ 87: 80], o60_10[ 79: 72], o60_11[ 79: 72], o60_12[ 79: 72], o60_13[ 79: 72],	o60_10[ 71: 64], o60_11[ 71: 64], o60_12[ 71: 64], o60_13[ 71: 64] };
		i60_22 <= { o60_10[ 63: 56], o60_11[ 63: 56], o60_12[ 63: 56], o60_13[ 63: 56], o60_10[ 55: 48], o60_11[ 55: 48], o60_12[ 55: 48], o60_13[ 55: 48], o60_10[ 47: 40], o60_11[ 47: 40], o60_12[ 47: 40], o60_13[ 47: 40], o60_10[ 39: 32], o60_11[ 39: 32], o60_12[ 39: 32], o60_13[ 39: 32] };
		i60_23 <= { o60_10[ 31: 24], o60_11[ 31: 24], o60_12[ 31: 24], o60_13[ 31: 24], o60_10[ 23: 16], o60_11[ 23: 16], o60_12[ 23: 16], o60_13[ 23: 16], o60_10[ 15:  8], o60_11[ 15:  8], o60_12[ 15:  8], o60_13[ 15:  8], o60_10[  7:  0], o60_11[  7:  0], o60_12[  7:  0], o60_13[  7:  0] };
		
	end

	reg  [127:0] i61_00, i61_01, i61_02, i61_03, i61_10, i61_11, i61_12, i61_13, i61_20, i61_21, i61_22, i61_23;
	wire [127:0] o61_00, o61_01, o61_02, o61_03, o61_10, o61_11, o61_12, o61_13, o61_20, o61_21, o61_22, o61_23;

	aes_round r61_00 (clk, i61_00, o61_00);
	aes_round r61_01 (clk, i61_01, o61_01);
	aes_round r61_02 (clk, i61_02, o61_02);
	aes_round r61_03 (clk, i61_03, o61_03);

	aes_round r61_10 (clk, i61_10, o61_10);
	aes_round r61_11 (clk, i61_11, o61_11);
	aes_round r61_12 (clk, i61_12, o61_12);
	aes_round r61_13 (clk, i61_13, o61_13);
	
	echo_mix  r61_20 (clk, i61_20, o61_20);
	echo_mix  r61_21 (clk, i61_21, o61_21);
	echo_mix  r61_22 (clk, i61_22, o61_22);
	echo_mix  r61_23 (clk, i61_23, o61_23);

	always @ ( posedge clk ) begin

		i61_00 <= { o51_20[127:120], o51_20[95:88], o51_20[63:56], o51_20[31:24], o51_21[127:120], o51_21[95:88], o51_21[63:56], o51_21[31:24], o51_22[127:120], o51_22[95:88], o51_22[63:56], o51_22[31:24], o51_23[127:120], o51_23[95:88], o51_23[63:56], o51_23[31:24] };
		i61_01 <= { o52_20[119:112], o52_20[87:80], o52_20[55:48], o52_20[23:16], o52_21[119:112], o52_21[87:80], o52_21[55:48], o52_21[23:16], o52_22[119:112], o52_22[87:80], o52_22[55:48], o52_22[23:16], o52_23[119:112], o52_23[87:80], o52_23[55:48], o52_23[23:16] };
		i61_02 <= { o53_20[111:104], o53_20[79:72], o53_20[47:40], o53_20[15: 8], o53_21[111:104], o53_21[79:72], o53_21[47:40], o53_21[15: 8], o53_22[111:104], o53_22[79:72], o53_22[47:40], o53_22[15: 8], o53_23[111:104], o53_23[79:72], o53_23[47:40], o53_23[15: 8] };
		i61_03 <= { o50_20[103: 96], o50_20[71:64], o50_20[39:32], o50_20[ 7: 0], o50_21[103: 96], o50_21[71:64], o50_21[39:32], o50_21[ 7: 0], o50_22[103: 96], o50_22[71:64], o50_22[39:32], o50_22[ 7: 0], o50_23[103: 96], o50_23[71:64], o50_23[39:32], o50_23[ 7: 0] };

		i61_10 <= { o61_00[127:108], o61_00[107:96] ^ 12'h0264, o61_00[95:0] };
		i61_11 <= { o61_01[127:108], o61_01[107:96] ^ 12'h0269, o61_01[95:0] };
		i61_12 <= { o61_02[127:108], o61_02[107:96] ^ 12'h026E, o61_02[95:0] };
		i61_13 <= { o61_03[127:108], o61_03[107:96] ^ 12'h0263, o61_03[95:0] };

		i61_20 <= { o61_10[127:120], o61_11[127:120], o61_12[127:120], o61_13[127:120], o61_10[119:112], o61_11[119:112], o61_12[119:112], o61_13[119:112], o61_10[111:104], o61_11[111:104], o61_12[111:104], o61_13[111:104], o61_10[103: 96], o61_11[103: 96], o61_12[103: 96], o61_13[103: 96] };
		i61_21 <= { o61_10[ 95: 88], o61_11[ 95: 88], o61_12[ 95: 88], o61_13[ 95: 88], o61_10[ 87: 80], o61_11[ 87: 80], o61_12[ 87: 80], o61_13[ 87: 80], o61_10[ 79: 72], o61_11[ 79: 72], o61_12[ 79: 72], o61_13[ 79: 72],	o61_10[ 71: 64], o61_11[ 71: 64], o61_12[ 71: 64], o61_13[ 71: 64] };
		i61_22 <= { o61_10[ 63: 56], o61_11[ 63: 56], o61_12[ 63: 56], o61_13[ 63: 56], o61_10[ 55: 48], o61_11[ 55: 48], o61_12[ 55: 48], o61_13[ 55: 48], o61_10[ 47: 40], o61_11[ 47: 40], o61_12[ 47: 40], o61_13[ 47: 40], o61_10[ 39: 32], o61_11[ 39: 32], o61_12[ 39: 32], o61_13[ 39: 32] };
		i61_23 <= { o61_10[ 31: 24], o61_11[ 31: 24], o61_12[ 31: 24], o61_13[ 31: 24], o61_10[ 23: 16], o61_11[ 23: 16], o61_12[ 23: 16], o61_13[ 23: 16], o61_10[ 15:  8], o61_11[ 15:  8], o61_12[ 15:  8], o61_13[ 15:  8], o61_10[  7:  0], o61_11[  7:  0], o61_12[  7:  0], o61_13[  7:  0] };

	end

	reg  [127:0] i62_00, i62_01, i62_02, i62_03, i62_10, i62_11, i62_12, i62_13, i62_20, i62_21, i62_22, i62_23;
	wire [127:0] o62_00, o62_01, o62_02, o62_03, o62_10, o62_11, o62_12, o62_13, o62_20, o62_21, o62_22, o62_23;

	aes_round r62_00 (clk, i62_00, o62_00);
	aes_round r62_01 (clk, i62_01, o62_01);
	aes_round r62_02 (clk, i62_02, o62_02);
	aes_round r62_03 (clk, i62_03, o62_03);

	aes_round r62_10 (clk, i62_10, o62_10);
	aes_round r62_11 (clk, i62_11, o62_11);
	aes_round r62_12 (clk, i62_12, o62_12);
	aes_round r62_13 (clk, i62_13, o62_13);
	
	echo_mix  r62_20 (clk, i62_20, o62_20);
	echo_mix  r62_21 (clk, i62_21, o62_21);
	echo_mix  r62_22 (clk, i62_22, o62_22);
	echo_mix  r62_23 (clk, i62_23, o62_23);

	always @ ( posedge clk ) begin

		i62_00 <= { o52_20[127:120], o52_20[95:88], o52_20[63:56], o52_20[31:24], o52_21[127:120], o52_21[95:88], o52_21[63:56], o52_21[31:24], o52_22[127:120], o52_22[95:88], o52_22[63:56], o52_22[31:24], o52_23[127:120], o52_23[95:88], o52_23[63:56], o52_23[31:24] };
		i62_01 <= { o53_20[119:112], o53_20[87:80], o53_20[55:48], o53_20[23:16], o53_21[119:112], o53_21[87:80], o53_21[55:48], o53_21[23:16], o53_22[119:112], o53_22[87:80], o53_22[55:48], o53_22[23:16], o53_23[119:112], o53_23[87:80], o53_23[55:48], o53_23[23:16] };
		i62_02 <= { o50_20[111:104], o50_20[79:72], o50_20[47:40], o50_20[15: 8], o50_21[111:104], o50_21[79:72], o50_21[47:40], o50_21[15: 8], o50_22[111:104], o50_22[79:72], o50_22[47:40], o50_22[15: 8], o50_23[111:104], o50_23[79:72], o50_23[47:40], o50_23[15: 8] };
		i62_03 <= { o51_20[103: 96], o51_20[71:64], o51_20[39:32], o51_20[ 7: 0], o51_21[103: 96], o51_21[71:64], o51_21[39:32], o51_21[ 7: 0], o51_22[103: 96], o51_22[71:64], o51_22[39:32], o51_22[ 7: 0], o51_23[103: 96], o51_23[71:64], o51_23[39:32], o51_23[ 7: 0] }; 

		i62_10 <= { o62_00[127:108], o62_00[107:96] ^ 12'h0268, o62_00[95:0] };
		i62_11 <= { o62_01[127:108], o62_01[107:96] ^ 12'h026D, o62_01[95:0] };
		i62_12 <= { o62_02[127:108], o62_02[107:96] ^ 12'h0262, o62_02[95:0] };
		i62_13 <= { o62_03[127:108], o62_03[107:96] ^ 12'h0267, o62_03[95:0] };

		i62_20 <= { o62_10[127:120], o62_11[127:120], o62_12[127:120], o62_13[127:120], o62_10[119:112], o62_11[119:112], o62_12[119:112], o62_13[119:112], o62_10[111:104], o62_11[111:104], o62_12[111:104], o62_13[111:104], o62_10[103: 96], o62_11[103: 96], o62_12[103: 96], o62_13[103: 96] };
		i62_21 <= { o62_10[ 95: 88], o62_11[ 95: 88], o62_12[ 95: 88], o62_13[ 95: 88], o62_10[ 87: 80], o62_11[ 87: 80], o62_12[ 87: 80], o62_13[ 87: 80], o62_10[ 79: 72], o62_11[ 79: 72], o62_12[ 79: 72], o62_13[ 79: 72],	o62_10[ 71: 64], o62_11[ 71: 64], o62_12[ 71: 64], o62_13[ 71: 64] };
		i62_22 <= { o62_10[ 63: 56], o62_11[ 63: 56], o62_12[ 63: 56], o62_13[ 63: 56], o62_10[ 55: 48], o62_11[ 55: 48], o62_12[ 55: 48], o62_13[ 55: 48], o62_10[ 47: 40], o62_11[ 47: 40], o62_12[ 47: 40], o62_13[ 47: 40], o62_10[ 39: 32], o62_11[ 39: 32], o62_12[ 39: 32], o62_13[ 39: 32] };
		i62_23 <= { o62_10[ 31: 24], o62_11[ 31: 24], o62_12[ 31: 24], o62_13[ 31: 24], o62_10[ 23: 16], o62_11[ 23: 16], o62_12[ 23: 16], o62_13[ 23: 16], o62_10[ 15:  8], o62_11[ 15:  8], o62_12[ 15:  8], o62_13[ 15:  8], o62_10[  7:  0], o62_11[  7:  0], o62_12[  7:  0], o62_13[  7:  0] };

	end

	reg  [127:0] i63_00, i63_01, i63_02, i63_03, i63_10, i63_11, i63_12, i63_13, i63_20, i63_21, i63_22, i63_23;
	wire [127:0] o63_00, o63_01, o63_02, o63_03, o63_10, o63_11, o63_12, o63_13, o63_20, o63_21, o63_22, o63_23;

	aes_round r63_00 (clk, i63_00, o63_00);
	aes_round r63_01 (clk, i63_01, o63_01);
	aes_round r63_02 (clk, i63_02, o63_02);
	aes_round r63_03 (clk, i63_03, o63_03);

	aes_round r63_10 (clk, i63_10, o63_10);
	aes_round r63_11 (clk, i63_11, o63_11);
	aes_round r63_12 (clk, i63_12, o63_12);
	aes_round r63_13 (clk, i63_13, o63_13);
	
	echo_mix  r63_20 (clk, i63_20, o63_20);
	echo_mix  r63_21 (clk, i63_21, o63_21);
	echo_mix  r63_22 (clk, i63_22, o63_22);
	echo_mix  r63_23 (clk, i63_23, o63_23);

	always @ ( posedge clk ) begin

		i63_00 <= { o53_20[127:120], o53_20[95:88], o53_20[63:56], o53_20[31:24], o53_21[127:120], o53_21[95:88], o53_21[63:56], o53_21[31:24], o53_22[127:120], o53_22[95:88], o53_22[63:56], o53_22[31:24], o53_23[127:120], o53_23[95:88], o53_23[63:56], o53_23[31:24] };
		i63_01 <= { o50_20[119:112], o50_20[87:80], o50_20[55:48], o50_20[23:16], o50_21[119:112], o50_21[87:80], o50_21[55:48], o50_21[23:16], o50_22[119:112], o50_22[87:80], o50_22[55:48], o50_22[23:16], o50_23[119:112], o50_23[87:80], o50_23[55:48], o50_23[23:16] };
		i63_02 <= { o51_20[111:104], o51_20[79:72], o51_20[47:40], o51_20[15: 8], o51_21[111:104], o51_21[79:72], o51_21[47:40], o51_21[15: 8], o51_22[111:104], o51_22[79:72], o51_22[47:40], o51_22[15: 8], o51_23[111:104], o51_23[79:72], o51_23[47:40], o51_23[15: 8] };
		i63_03 <= { o52_20[103: 96], o52_20[71:64], o52_20[39:32], o52_20[ 7: 0], o52_21[103: 96], o52_21[71:64], o52_21[39:32], o52_21[ 7: 0], o52_22[103: 96], o52_22[71:64], o52_22[39:32], o52_22[ 7: 0], o52_23[103: 96], o52_23[71:64], o52_23[39:32], o52_23[ 7: 0] }; 

		i63_10 <= { o63_00[127:108], o63_00[107:96] ^ 12'h026C, o63_00[95:0] };
		i63_11 <= { o63_01[127:108], o63_01[107:96] ^ 12'h0261, o63_01[95:0] };
		i63_12 <= { o63_02[127:108], o63_02[107:96] ^ 12'h0266, o63_02[95:0] };
		i63_13 <= { o63_03[127:108], o63_03[107:96] ^ 12'h026B, o63_03[95:0] };

		i63_20 <= { o63_10[127:120], o63_11[127:120], o63_12[127:120], o63_13[127:120], o63_10[119:112], o63_11[119:112], o63_12[119:112], o63_13[119:112], o63_10[111:104], o63_11[111:104], o63_12[111:104], o63_13[111:104], o63_10[103: 96], o63_11[103: 96], o63_12[103: 96], o63_13[103: 96] };
		i63_21 <= { o63_10[ 95: 88], o63_11[ 95: 88], o63_12[ 95: 88], o63_13[ 95: 88], o63_10[ 87: 80], o63_11[ 87: 80], o63_12[ 87: 80], o63_13[ 87: 80], o63_10[ 79: 72], o63_11[ 79: 72], o63_12[ 79: 72], o63_13[ 79: 72],	o63_10[ 71: 64], o63_11[ 71: 64], o63_12[ 71: 64], o63_13[ 71: 64] };
		i63_22 <= { o63_10[ 63: 56], o63_11[ 63: 56], o63_12[ 63: 56], o63_13[ 63: 56], o63_10[ 55: 48], o63_11[ 55: 48], o63_12[ 55: 48], o63_13[ 55: 48], o63_10[ 47: 40], o63_11[ 47: 40], o63_12[ 47: 40], o63_13[ 47: 40], o63_10[ 39: 32], o63_11[ 39: 32], o63_12[ 39: 32], o63_13[ 39: 32] };
		i63_23 <= { o63_10[ 31: 24], o63_11[ 31: 24], o63_12[ 31: 24], o63_13[ 31: 24], o63_10[ 23: 16], o63_11[ 23: 16], o63_12[ 23: 16], o63_13[ 23: 16], o63_10[ 15:  8], o63_11[ 15:  8], o63_12[ 15:  8], o63_13[ 15:  8], o63_10[  7:  0], o63_11[  7:  0], o63_12[  7:  0], o63_13[  7:  0] };

	end

	// ROUND 7

	reg  [127:0] i70_00, i70_01, i70_02, i70_03, i70_10, i70_11, i70_12, i70_13, i70_20, i70_21, i70_22, i70_23;
	wire [127:0] o70_00, o70_01, o70_02, o70_03, o70_10, o70_11, o70_12, o70_13, o70_20, o70_21, o70_22, o70_23;

	aes_round r70_00 (clk, i70_00, o70_00);
	aes_round r70_01 (clk, i70_01, o70_01);
	aes_round r70_02 (clk, i70_02, o70_02);
	aes_round r70_03 (clk, i70_03, o70_03);

	aes_round r70_10 (clk, i70_10, o70_10);
	aes_round r70_11 (clk, i70_11, o70_11);
	aes_round r70_12 (clk, i70_12, o70_12);
	aes_round r70_13 (clk, i70_13, o70_13);
	
	echo_mix  r70_20 (clk, i70_20, o70_20);
	echo_mix  r70_21 (clk, i70_21, o70_21);
	echo_mix  r70_22 (clk, i70_22, o70_22);
	echo_mix  r70_23 (clk, i70_23, o70_23);

	always @ ( posedge clk ) begin

		i70_00 <= { o60_20[127:120], o60_20[95:88], o60_20[63:56], o60_20[31:24], o60_21[127:120], o60_21[95:88], o60_21[63:56], o60_21[31:24], o60_22[127:120], o60_22[95:88], o60_22[63:56], o60_22[31:24], o60_23[127:120], o60_23[95:88], o60_23[63:56], o60_23[31:24] };
		i70_01 <= { o61_20[119:112], o61_20[87:80], o61_20[55:48], o61_20[23:16], o61_21[119:112], o61_21[87:80], o61_21[55:48], o61_21[23:16], o61_22[119:112], o61_22[87:80], o61_22[55:48], o61_22[23:16], o61_23[119:112], o61_23[87:80], o61_23[55:48], o61_23[23:16] };
		i70_02 <= { o62_20[111:104], o62_20[79:72], o62_20[47:40], o62_20[15: 8], o62_21[111:104], o62_21[79:72], o62_21[47:40], o62_21[15: 8], o62_22[111:104], o62_22[79:72], o62_22[47:40], o62_22[15: 8], o62_23[111:104], o62_23[79:72], o62_23[47:40], o62_23[15: 8] };
		i70_03 <= { o63_20[103: 96], o63_20[71:64], o63_20[39:32], o63_20[ 7: 0], o63_21[103: 96], o63_21[71:64], o63_21[39:32], o63_21[ 7: 0], o63_22[103: 96], o63_22[71:64], o63_22[39:32], o63_22[ 7: 0], o63_23[103: 96], o63_23[71:64], o63_23[39:32], o63_23[ 7: 0] }; 

		i70_10 <= { o70_00[127:108], o70_00[107:96] ^ 12'h0270, o70_00[95:0] };
		i70_11 <= { o70_01[127:108], o70_01[107:96] ^ 12'h0275, o70_01[95:0] };
		i70_12 <= { o70_02[127:108], o70_02[107:96] ^ 12'h027A, o70_02[95:0] };
		i70_13 <= { o70_03[127:108], o70_03[107:96] ^ 12'h027F, o70_03[95:0] };

		i70_20 <= { o70_10[127:120], o70_11[127:120], o70_12[127:120], o70_13[127:120], o70_10[119:112], o70_11[119:112], o70_12[119:112], o70_13[119:112], o70_10[111:104], o70_11[111:104], o70_12[111:104], o70_13[111:104], o70_10[103: 96], o70_11[103: 96], o70_12[103: 96], o70_13[103: 96] };
		i70_21 <= { o70_10[ 95: 88], o70_11[ 95: 88], o70_12[ 95: 88], o70_13[ 95: 88], o70_10[ 87: 80], o70_11[ 87: 80], o70_12[ 87: 80], o70_13[ 87: 80], o70_10[ 79: 72], o70_11[ 79: 72], o70_12[ 79: 72], o70_13[ 79: 72],	o70_10[ 71: 64], o70_11[ 71: 64], o70_12[ 71: 64], o70_13[ 71: 64] };
		i70_22 <= { o70_10[ 63: 56], o70_11[ 63: 56], o70_12[ 63: 56], o70_13[ 63: 56], o70_10[ 55: 48], o70_11[ 55: 48], o70_12[ 55: 48], o70_13[ 55: 48], o70_10[ 47: 40], o70_11[ 47: 40], o70_12[ 47: 40], o70_13[ 47: 40], o70_10[ 39: 32], o70_11[ 39: 32], o70_12[ 39: 32], o70_13[ 39: 32] };
		i70_23 <= { o70_10[ 31: 24], o70_11[ 31: 24], o70_12[ 31: 24], o70_13[ 31: 24], o70_10[ 23: 16], o70_11[ 23: 16], o70_12[ 23: 16], o70_13[ 23: 16], o70_10[ 15:  8], o70_11[ 15:  8], o70_12[ 15:  8], o70_13[ 15:  8], o70_10[  7:  0], o70_11[  7:  0], o70_12[  7:  0], o70_13[  7:  0] };
		
	end

	reg  [127:0] i71_00, i71_01, i71_02, i71_03, i71_10, i71_11, i71_12, i71_13, i71_20, i71_21, i71_22, i71_23;
	wire [127:0] o71_00, o71_01, o71_02, o71_03, o71_10, o71_11, o71_12, o71_13, o71_20, o71_21, o71_22, o71_23;

	aes_round r71_00 (clk, i71_00, o71_00);
	aes_round r71_01 (clk, i71_01, o71_01);
	aes_round r71_02 (clk, i71_02, o71_02);
	aes_round r71_03 (clk, i71_03, o71_03);

	aes_round r71_10 (clk, i71_10, o71_10);
	aes_round r71_11 (clk, i71_11, o71_11);
	aes_round r71_12 (clk, i71_12, o71_12);
	aes_round r71_13 (clk, i71_13, o71_13);
	
	echo_mix  r71_20 (clk, i71_20, o71_20);
	echo_mix  r71_21 (clk, i71_21, o71_21);
	echo_mix  r71_22 (clk, i71_22, o71_22);
	echo_mix  r71_23 (clk, i71_23, o71_23);

	always @ ( posedge clk ) begin

		i71_00 <= { o61_20[127:120], o61_20[95:88], o61_20[63:56], o61_20[31:24], o61_21[127:120], o61_21[95:88], o61_21[63:56], o61_21[31:24], o61_22[127:120], o61_22[95:88], o61_22[63:56], o61_22[31:24], o61_23[127:120], o61_23[95:88], o61_23[63:56], o61_23[31:24] };
		i71_01 <= { o62_20[119:112], o62_20[87:80], o62_20[55:48], o62_20[23:16], o62_21[119:112], o62_21[87:80], o62_21[55:48], o62_21[23:16], o62_22[119:112], o62_22[87:80], o62_22[55:48], o62_22[23:16], o62_23[119:112], o62_23[87:80], o62_23[55:48], o62_23[23:16] };
		i71_02 <= { o63_20[111:104], o63_20[79:72], o63_20[47:40], o63_20[15: 8], o63_21[111:104], o63_21[79:72], o63_21[47:40], o63_21[15: 8], o63_22[111:104], o63_22[79:72], o63_22[47:40], o63_22[15: 8], o63_23[111:104], o63_23[79:72], o63_23[47:40], o63_23[15: 8] };
		i71_03 <= { o60_20[103: 96], o60_20[71:64], o60_20[39:32], o60_20[ 7: 0], o60_21[103: 96], o60_21[71:64], o60_21[39:32], o60_21[ 7: 0], o60_22[103: 96], o60_22[71:64], o60_22[39:32], o60_22[ 7: 0], o60_23[103: 96], o60_23[71:64], o60_23[39:32], o60_23[ 7: 0] };

		i71_10 <= { o71_00[127:108], o71_00[107:96] ^ 12'h0274, o71_00[95:0] };
		i71_11 <= { o71_01[127:108], o71_01[107:96] ^ 12'h0279, o71_01[95:0] };
		i71_12 <= { o71_02[127:108], o71_02[107:96] ^ 12'h027E, o71_02[95:0] };
		i71_13 <= { o71_03[127:108], o71_03[107:96] ^ 12'h0273, o71_03[95:0] };

		i71_20 <= { o71_10[127:120], o71_11[127:120], o71_12[127:120], o71_13[127:120], o71_10[119:112], o71_11[119:112], o71_12[119:112], o71_13[119:112], o71_10[111:104], o71_11[111:104], o71_12[111:104], o71_13[111:104], o71_10[103: 96], o71_11[103: 96], o71_12[103: 96], o71_13[103: 96] };
		i71_21 <= { o71_10[ 95: 88], o71_11[ 95: 88], o71_12[ 95: 88], o71_13[ 95: 88], o71_10[ 87: 80], o71_11[ 87: 80], o71_12[ 87: 80], o71_13[ 87: 80], o71_10[ 79: 72], o71_11[ 79: 72], o71_12[ 79: 72], o71_13[ 79: 72],	o71_10[ 71: 64], o71_11[ 71: 64], o71_12[ 71: 64], o71_13[ 71: 64] };
		i71_22 <= { o71_10[ 63: 56], o71_11[ 63: 56], o71_12[ 63: 56], o71_13[ 63: 56], o71_10[ 55: 48], o71_11[ 55: 48], o71_12[ 55: 48], o71_13[ 55: 48], o71_10[ 47: 40], o71_11[ 47: 40], o71_12[ 47: 40], o71_13[ 47: 40], o71_10[ 39: 32], o71_11[ 39: 32], o71_12[ 39: 32], o71_13[ 39: 32] };
		i71_23 <= { o71_10[ 31: 24], o71_11[ 31: 24], o71_12[ 31: 24], o71_13[ 31: 24], o71_10[ 23: 16], o71_11[ 23: 16], o71_12[ 23: 16], o71_13[ 23: 16], o71_10[ 15:  8], o71_11[ 15:  8], o71_12[ 15:  8], o71_13[ 15:  8], o71_10[  7:  0], o71_11[  7:  0], o71_12[  7:  0], o71_13[  7:  0] };

	end

	reg  [127:0] i72_00, i72_01, i72_02, i72_03, i72_10, i72_11, i72_12, i72_13, i72_20, i72_21, i72_22, i72_23;
	wire [127:0] o72_00, o72_01, o72_02, o72_03, o72_10, o72_11, o72_12, o72_13, o72_20, o72_21, o72_22, o72_23;

	aes_round r72_00 (clk, i72_00, o72_00);
	aes_round r72_01 (clk, i72_01, o72_01);
	aes_round r72_02 (clk, i72_02, o72_02);
	aes_round r72_03 (clk, i72_03, o72_03);

	aes_round r72_10 (clk, i72_10, o72_10);
	aes_round r72_11 (clk, i72_11, o72_11);
	aes_round r72_12 (clk, i72_12, o72_12);
	aes_round r72_13 (clk, i72_13, o72_13);
	
	echo_mix  r72_20 (clk, i72_20, o72_20);
	echo_mix  r72_21 (clk, i72_21, o72_21);
	echo_mix  r72_22 (clk, i72_22, o72_22);
	echo_mix  r72_23 (clk, i72_23, o72_23);

	always @ ( posedge clk ) begin

		i72_00 <= { o62_20[127:120], o62_20[95:88], o62_20[63:56], o62_20[31:24], o62_21[127:120], o62_21[95:88], o62_21[63:56], o62_21[31:24], o62_22[127:120], o62_22[95:88], o62_22[63:56], o62_22[31:24], o62_23[127:120], o62_23[95:88], o62_23[63:56], o62_23[31:24] };
		i72_01 <= { o63_20[119:112], o63_20[87:80], o63_20[55:48], o63_20[23:16], o63_21[119:112], o63_21[87:80], o63_21[55:48], o63_21[23:16], o63_22[119:112], o63_22[87:80], o63_22[55:48], o63_22[23:16], o63_23[119:112], o63_23[87:80], o63_23[55:48], o63_23[23:16] };
		i72_02 <= { o60_20[111:104], o60_20[79:72], o60_20[47:40], o60_20[15: 8], o60_21[111:104], o60_21[79:72], o60_21[47:40], o60_21[15: 8], o60_22[111:104], o60_22[79:72], o60_22[47:40], o60_22[15: 8], o60_23[111:104], o60_23[79:72], o60_23[47:40], o60_23[15: 8] };
		i72_03 <= { o61_20[103: 96], o61_20[71:64], o61_20[39:32], o61_20[ 7: 0], o61_21[103: 96], o61_21[71:64], o61_21[39:32], o61_21[ 7: 0], o61_22[103: 96], o61_22[71:64], o61_22[39:32], o61_22[ 7: 0], o61_23[103: 96], o61_23[71:64], o61_23[39:32], o61_23[ 7: 0] }; 

		i72_10 <= { o72_00[127:108], o72_00[107:96] ^ 12'h0278, o72_00[95:0] };
		i72_11 <= { o72_01[127:108], o72_01[107:96] ^ 12'h027D, o72_01[95:0] };
		i72_12 <= { o72_02[127:108], o72_02[107:96] ^ 12'h0272, o72_02[95:0] };
		i72_13 <= { o72_03[127:108], o72_03[107:96] ^ 12'h0277, o72_03[95:0] };

		i72_20 <= { o72_10[127:120], o72_11[127:120], o72_12[127:120], o72_13[127:120], o72_10[119:112], o72_11[119:112], o72_12[119:112], o72_13[119:112], o72_10[111:104], o72_11[111:104], o72_12[111:104], o72_13[111:104], o72_10[103: 96], o72_11[103: 96], o72_12[103: 96], o72_13[103: 96] };
		i72_21 <= { o72_10[ 95: 88], o72_11[ 95: 88], o72_12[ 95: 88], o72_13[ 95: 88], o72_10[ 87: 80], o72_11[ 87: 80], o72_12[ 87: 80], o72_13[ 87: 80], o72_10[ 79: 72], o72_11[ 79: 72], o72_12[ 79: 72], o72_13[ 79: 72],	o72_10[ 71: 64], o72_11[ 71: 64], o72_12[ 71: 64], o72_13[ 71: 64] };
		i72_22 <= { o72_10[ 63: 56], o72_11[ 63: 56], o72_12[ 63: 56], o72_13[ 63: 56], o72_10[ 55: 48], o72_11[ 55: 48], o72_12[ 55: 48], o72_13[ 55: 48], o72_10[ 47: 40], o72_11[ 47: 40], o72_12[ 47: 40], o72_13[ 47: 40], o72_10[ 39: 32], o72_11[ 39: 32], o72_12[ 39: 32], o72_13[ 39: 32] };
		i72_23 <= { o72_10[ 31: 24], o72_11[ 31: 24], o72_12[ 31: 24], o72_13[ 31: 24], o72_10[ 23: 16], o72_11[ 23: 16], o72_12[ 23: 16], o72_13[ 23: 16], o72_10[ 15:  8], o72_11[ 15:  8], o72_12[ 15:  8], o72_13[ 15:  8], o72_10[  7:  0], o72_11[  7:  0], o72_12[  7:  0], o72_13[  7:  0] };

	end

	reg  [127:0] i73_00, i73_01, i73_02, i73_03, i73_10, i73_11, i73_12, i73_13, i73_20, i73_21, i73_22, i73_23;
	wire [127:0] o73_00, o73_01, o73_02, o73_03, o73_10, o73_11, o73_12, o73_13, o73_20, o73_21, o73_22, o73_23;

	aes_round r73_00 (clk, i73_00, o73_00);
	aes_round r73_01 (clk, i73_01, o73_01);
	aes_round r73_02 (clk, i73_02, o73_02);
	aes_round r73_03 (clk, i73_03, o73_03);

	aes_round r73_10 (clk, i73_10, o73_10);
	aes_round r73_11 (clk, i73_11, o73_11);
	aes_round r73_12 (clk, i73_12, o73_12);
	aes_round r73_13 (clk, i73_13, o73_13);
	
	echo_mix  r73_20 (clk, i73_20, o73_20);
	echo_mix  r73_21 (clk, i73_21, o73_21);
	echo_mix  r73_22 (clk, i73_22, o73_22);
	echo_mix  r73_23 (clk, i73_23, o73_23);

	always @ ( posedge clk ) begin

		i73_00 <= { o63_20[127:120], o63_20[95:88], o63_20[63:56], o63_20[31:24], o63_21[127:120], o63_21[95:88], o63_21[63:56], o63_21[31:24], o63_22[127:120], o63_22[95:88], o63_22[63:56], o63_22[31:24], o63_23[127:120], o63_23[95:88], o63_23[63:56], o63_23[31:24] };
		i73_01 <= { o60_20[119:112], o60_20[87:80], o60_20[55:48], o60_20[23:16], o60_21[119:112], o60_21[87:80], o60_21[55:48], o60_21[23:16], o60_22[119:112], o60_22[87:80], o60_22[55:48], o60_22[23:16], o60_23[119:112], o60_23[87:80], o60_23[55:48], o60_23[23:16] };
		i73_02 <= { o61_20[111:104], o61_20[79:72], o61_20[47:40], o61_20[15: 8], o61_21[111:104], o61_21[79:72], o61_21[47:40], o61_21[15: 8], o61_22[111:104], o61_22[79:72], o61_22[47:40], o61_22[15: 8], o61_23[111:104], o61_23[79:72], o61_23[47:40], o61_23[15: 8] };
		i73_03 <= { o62_20[103: 96], o62_20[71:64], o62_20[39:32], o62_20[ 7: 0], o62_21[103: 96], o62_21[71:64], o62_21[39:32], o62_21[ 7: 0], o62_22[103: 96], o62_22[71:64], o62_22[39:32], o62_22[ 7: 0], o62_23[103: 96], o62_23[71:64], o62_23[39:32], o62_23[ 7: 0] }; 

		i73_10 <= { o73_00[127:108], o73_00[107:96] ^ 12'h027C, o73_00[95:0] };
		i73_11 <= { o73_01[127:108], o73_01[107:96] ^ 12'h0271, o73_01[95:0] };
		i73_12 <= { o73_02[127:108], o73_02[107:96] ^ 12'h0276, o73_02[95:0] };
		i73_13 <= { o73_03[127:108], o73_03[107:96] ^ 12'h027B, o73_03[95:0] };

		i73_20 <= { o73_10[127:120], o73_11[127:120], o73_12[127:120], o73_13[127:120], o73_10[119:112], o73_11[119:112], o73_12[119:112], o73_13[119:112], o73_10[111:104], o73_11[111:104], o73_12[111:104], o73_13[111:104], o73_10[103: 96], o73_11[103: 96], o73_12[103: 96], o73_13[103: 96] };
		i73_21 <= { o73_10[ 95: 88], o73_11[ 95: 88], o73_12[ 95: 88], o73_13[ 95: 88], o73_10[ 87: 80], o73_11[ 87: 80], o73_12[ 87: 80], o73_13[ 87: 80], o73_10[ 79: 72], o73_11[ 79: 72], o73_12[ 79: 72], o73_13[ 79: 72],	o73_10[ 71: 64], o73_11[ 71: 64], o73_12[ 71: 64], o73_13[ 71: 64] };
		i73_22 <= { o73_10[ 63: 56], o73_11[ 63: 56], o73_12[ 63: 56], o73_13[ 63: 56], o73_10[ 55: 48], o73_11[ 55: 48], o73_12[ 55: 48], o73_13[ 55: 48], o73_10[ 47: 40], o73_11[ 47: 40], o73_12[ 47: 40], o73_13[ 47: 40], o73_10[ 39: 32], o73_11[ 39: 32], o73_12[ 39: 32], o73_13[ 39: 32] };
		i73_23 <= { o73_10[ 31: 24], o73_11[ 31: 24], o73_12[ 31: 24], o73_13[ 31: 24], o73_10[ 23: 16], o73_11[ 23: 16], o73_12[ 23: 16], o73_13[ 23: 16], o73_10[ 15:  8], o73_11[ 15:  8], o73_12[ 15:  8], o73_13[ 15:  8], o73_10[  7:  0], o73_11[  7:  0], o73_12[  7:  0], o73_13[  7:  0] };

	end

	// ROUND 8

	reg  [127:0] i80_00, i80_01, i80_02, i80_03, i80_10, i80_11, i80_12, i80_13, i80_20, i80_21, i80_22, i80_23;
	wire [127:0] o80_00, o80_01, o80_02, o80_03, o80_10, o80_11, o80_12, o80_13, o80_20, o80_21, o80_22, o80_23;

	aes_round r80_00 (clk, i80_00, o80_00);
	aes_round r80_01 (clk, i80_01, o80_01);
	aes_round r80_02 (clk, i80_02, o80_02);
	aes_round r80_03 (clk, i80_03, o80_03);

	aes_round r80_10 (clk, i80_10, o80_10);
	aes_round r80_11 (clk, i80_11, o80_11);
	aes_round r80_12 (clk, i80_12, o80_12);
	aes_round r80_13 (clk, i80_13, o80_13);
	
	echo_mix  r80_20 (clk, i80_20, o80_20);
	echo_mix  r80_21 (clk, i80_21, o80_21);
	echo_mix  r80_22 (clk, i80_22, o80_22);
	echo_mix  r80_23 (clk, i80_23, o80_23);

	always @ ( posedge clk ) begin

		i80_00 <= { o70_20[127:120], o70_20[95:88], o70_20[63:56], o70_20[31:24], o70_21[127:120], o70_21[95:88], o70_21[63:56], o70_21[31:24], o70_22[127:120], o70_22[95:88], o70_22[63:56], o70_22[31:24], o70_23[127:120], o70_23[95:88], o70_23[63:56], o70_23[31:24] };
		i80_01 <= { o71_20[119:112], o71_20[87:80], o71_20[55:48], o71_20[23:16], o71_21[119:112], o71_21[87:80], o71_21[55:48], o71_21[23:16], o71_22[119:112], o71_22[87:80], o71_22[55:48], o71_22[23:16], o71_23[119:112], o71_23[87:80], o71_23[55:48], o71_23[23:16] };
		i80_02 <= { o72_20[111:104], o72_20[79:72], o72_20[47:40], o72_20[15: 8], o72_21[111:104], o72_21[79:72], o72_21[47:40], o72_21[15: 8], o72_22[111:104], o72_22[79:72], o72_22[47:40], o72_22[15: 8], o72_23[111:104], o72_23[79:72], o72_23[47:40], o72_23[15: 8] };
		i80_03 <= { o73_20[103: 96], o73_20[71:64], o73_20[39:32], o73_20[ 7: 0], o73_21[103: 96], o73_21[71:64], o73_21[39:32], o73_21[ 7: 0], o73_22[103: 96], o73_22[71:64], o73_22[39:32], o73_22[ 7: 0], o73_23[103: 96], o73_23[71:64], o73_23[39:32], o73_23[ 7: 0] }; 

		i80_10 <= { o80_00[127:108], o80_00[107:96] ^ 12'h0280, o80_00[95:0] };
		i80_11 <= { o80_01[127:108], o80_01[107:96] ^ 12'h0285, o80_01[95:0] };
		i80_12 <= { o80_02[127:108], o80_02[107:96] ^ 12'h028A, o80_02[95:0] };
		i80_13 <= { o80_03[127:108], o80_03[107:96] ^ 12'h028F, o80_03[95:0] };

		i80_20 <= { o80_10[127:120], o80_11[127:120], o80_12[127:120], o80_13[127:120], o80_10[119:112], o80_11[119:112], o80_12[119:112], o80_13[119:112], o80_10[111:104], o80_11[111:104], o80_12[111:104], o80_13[111:104], o80_10[103: 96], o80_11[103: 96], o80_12[103: 96], o80_13[103: 96] };
		i80_21 <= { o80_10[ 95: 88], o80_11[ 95: 88], o80_12[ 95: 88], o80_13[ 95: 88], o80_10[ 87: 80], o80_11[ 87: 80], o80_12[ 87: 80], o80_13[ 87: 80], o80_10[ 79: 72], o80_11[ 79: 72], o80_12[ 79: 72], o80_13[ 79: 72],	o80_10[ 71: 64], o80_11[ 71: 64], o80_12[ 71: 64], o80_13[ 71: 64] };
		i80_22 <= { o80_10[ 63: 56], o80_11[ 63: 56], o80_12[ 63: 56], o80_13[ 63: 56], o80_10[ 55: 48], o80_11[ 55: 48], o80_12[ 55: 48], o80_13[ 55: 48], o80_10[ 47: 40], o80_11[ 47: 40], o80_12[ 47: 40], o80_13[ 47: 40], o80_10[ 39: 32], o80_11[ 39: 32], o80_12[ 39: 32], o80_13[ 39: 32] };
		i80_23 <= { o80_10[ 31: 24], o80_11[ 31: 24], o80_12[ 31: 24], o80_13[ 31: 24], o80_10[ 23: 16], o80_11[ 23: 16], o80_12[ 23: 16], o80_13[ 23: 16], o80_10[ 15:  8], o80_11[ 15:  8], o80_12[ 15:  8], o80_13[ 15:  8], o80_10[  7:  0], o80_11[  7:  0], o80_12[  7:  0], o80_13[  7:  0] };
		
	end

	reg  [127:0] i81_00, i81_01, i81_02, i81_03, i81_10, i81_11, i81_12, i81_13, i81_20, i81_21, i81_22, i81_23;
	wire [127:0] o81_00, o81_01, o81_02, o81_03, o81_10, o81_11, o81_12, o81_13, o81_20, o81_21, o81_22, o81_23;

	aes_round r81_00 (clk, i81_00, o81_00);
	aes_round r81_01 (clk, i81_01, o81_01);
	aes_round r81_02 (clk, i81_02, o81_02);
	aes_round r81_03 (clk, i81_03, o81_03);

	aes_round r81_10 (clk, i81_10, o81_10);
	aes_round r81_11 (clk, i81_11, o81_11);
	aes_round r81_12 (clk, i81_12, o81_12);
	aes_round r81_13 (clk, i81_13, o81_13);
	
	echo_mix  r81_20 (clk, i81_20, o81_20);
	echo_mix  r81_21 (clk, i81_21, o81_21);
	echo_mix  r81_22 (clk, i81_22, o81_22);
	echo_mix  r81_23 (clk, i81_23, o81_23);

	always @ ( posedge clk ) begin

		i81_00 <= { o71_20[127:120], o71_20[95:88], o71_20[63:56], o71_20[31:24], o71_21[127:120], o71_21[95:88], o71_21[63:56], o71_21[31:24], o71_22[127:120], o71_22[95:88], o71_22[63:56], o71_22[31:24], o71_23[127:120], o71_23[95:88], o71_23[63:56], o71_23[31:24] };
		i81_01 <= { o72_20[119:112], o72_20[87:80], o72_20[55:48], o72_20[23:16], o72_21[119:112], o72_21[87:80], o72_21[55:48], o72_21[23:16], o72_22[119:112], o72_22[87:80], o72_22[55:48], o72_22[23:16], o72_23[119:112], o72_23[87:80], o72_23[55:48], o72_23[23:16] };
		i81_02 <= { o73_20[111:104], o73_20[79:72], o73_20[47:40], o73_20[15: 8], o73_21[111:104], o73_21[79:72], o73_21[47:40], o73_21[15: 8], o73_22[111:104], o73_22[79:72], o73_22[47:40], o73_22[15: 8], o73_23[111:104], o73_23[79:72], o73_23[47:40], o73_23[15: 8] };
		i81_03 <= { o70_20[103: 96], o70_20[71:64], o70_20[39:32], o70_20[ 7: 0], o70_21[103: 96], o70_21[71:64], o70_21[39:32], o70_21[ 7: 0], o70_22[103: 96], o70_22[71:64], o70_22[39:32], o70_22[ 7: 0], o70_23[103: 96], o70_23[71:64], o70_23[39:32], o70_23[ 7: 0] };

		i81_10 <= { o81_00[127:108], o81_00[107:96] ^ 12'h0284, o81_00[95:0] };
		i81_11 <= { o81_01[127:108], o81_01[107:96] ^ 12'h0289, o81_01[95:0] };
		i81_12 <= { o81_02[127:108], o81_02[107:96] ^ 12'h028E, o81_02[95:0] };
		i81_13 <= { o81_03[127:108], o81_03[107:96] ^ 12'h0283, o81_03[95:0] };

		i81_20 <= { o81_10[127:120], o81_11[127:120], o81_12[127:120], o81_13[127:120], o81_10[119:112], o81_11[119:112], o81_12[119:112], o81_13[119:112], o81_10[111:104], o81_11[111:104], o81_12[111:104], o81_13[111:104], o81_10[103: 96], o81_11[103: 96], o81_12[103: 96], o81_13[103: 96] };
		i81_21 <= { o81_10[ 95: 88], o81_11[ 95: 88], o81_12[ 95: 88], o81_13[ 95: 88], o81_10[ 87: 80], o81_11[ 87: 80], o81_12[ 87: 80], o81_13[ 87: 80], o81_10[ 79: 72], o81_11[ 79: 72], o81_12[ 79: 72], o81_13[ 79: 72],	o81_10[ 71: 64], o81_11[ 71: 64], o81_12[ 71: 64], o81_13[ 71: 64] };
		i81_22 <= { o81_10[ 63: 56], o81_11[ 63: 56], o81_12[ 63: 56], o81_13[ 63: 56], o81_10[ 55: 48], o81_11[ 55: 48], o81_12[ 55: 48], o81_13[ 55: 48], o81_10[ 47: 40], o81_11[ 47: 40], o81_12[ 47: 40], o81_13[ 47: 40], o81_10[ 39: 32], o81_11[ 39: 32], o81_12[ 39: 32], o81_13[ 39: 32] };
		i81_23 <= { o81_10[ 31: 24], o81_11[ 31: 24], o81_12[ 31: 24], o81_13[ 31: 24], o81_10[ 23: 16], o81_11[ 23: 16], o81_12[ 23: 16], o81_13[ 23: 16], o81_10[ 15:  8], o81_11[ 15:  8], o81_12[ 15:  8], o81_13[ 15:  8], o81_10[  7:  0], o81_11[  7:  0], o81_12[  7:  0], o81_13[  7:  0] };

	end

	reg  [127:0] i82_00, i82_01, i82_02, i82_03, i82_10, i82_11, i82_12, i82_13, i82_20, i82_21, i82_22, i82_23;
	wire [127:0] o82_00, o82_01, o82_02, o82_03, o82_10, o82_11, o82_12, o82_13, o82_20, o82_21, o82_22, o82_23;

	aes_round r82_00 (clk, i82_00, o82_00);
	aes_round r82_01 (clk, i82_01, o82_01);
	aes_round r82_02 (clk, i82_02, o82_02);
	aes_round r82_03 (clk, i82_03, o82_03);

	aes_round r82_10 (clk, i82_10, o82_10);
	aes_round r82_11 (clk, i82_11, o82_11);
	aes_round r82_12 (clk, i82_12, o82_12);
	aes_round r82_13 (clk, i82_13, o82_13);
	
	echo_mix  r82_20 (clk, i82_20, o82_20);
	echo_mix  r82_21 (clk, i82_21, o82_21);
	echo_mix  r82_22 (clk, i82_22, o82_22);
	echo_mix  r82_23 (clk, i82_23, o82_23);

	always @ ( posedge clk ) begin

		i82_00 <= { o72_20[127:120], o72_20[95:88], o72_20[63:56], o72_20[31:24], o72_21[127:120], o72_21[95:88], o72_21[63:56], o72_21[31:24], o72_22[127:120], o72_22[95:88], o72_22[63:56], o72_22[31:24], o72_23[127:120], o72_23[95:88], o72_23[63:56], o72_23[31:24] };
		i82_01 <= { o73_20[119:112], o73_20[87:80], o73_20[55:48], o73_20[23:16], o73_21[119:112], o73_21[87:80], o73_21[55:48], o73_21[23:16], o73_22[119:112], o73_22[87:80], o73_22[55:48], o73_22[23:16], o73_23[119:112], o73_23[87:80], o73_23[55:48], o73_23[23:16] };
		i82_02 <= { o70_20[111:104], o70_20[79:72], o70_20[47:40], o70_20[15: 8], o70_21[111:104], o70_21[79:72], o70_21[47:40], o70_21[15: 8], o70_22[111:104], o70_22[79:72], o70_22[47:40], o70_22[15: 8], o70_23[111:104], o70_23[79:72], o70_23[47:40], o70_23[15: 8] };
		i82_03 <= { o71_20[103: 96], o71_20[71:64], o71_20[39:32], o71_20[ 7: 0], o71_21[103: 96], o71_21[71:64], o71_21[39:32], o71_21[ 7: 0], o71_22[103: 96], o71_22[71:64], o71_22[39:32], o71_22[ 7: 0], o71_23[103: 96], o71_23[71:64], o71_23[39:32], o71_23[ 7: 0] }; 

		i82_10 <= { o82_00[127:108], o82_00[107:96] ^ 12'h0288, o82_00[95:0] };
		i82_11 <= { o82_01[127:108], o82_01[107:96] ^ 12'h028D, o82_01[95:0] };
		i82_12 <= { o82_02[127:108], o82_02[107:96] ^ 12'h0282, o82_02[95:0] };
		i82_13 <= { o82_03[127:108], o82_03[107:96] ^ 12'h0287, o82_03[95:0] };

		i82_20 <= { o82_10[127:120], o82_11[127:120], o82_12[127:120], o82_13[127:120], o82_10[119:112], o82_11[119:112], o82_12[119:112], o82_13[119:112], o82_10[111:104], o82_11[111:104], o82_12[111:104], o82_13[111:104], o82_10[103: 96], o82_11[103: 96], o82_12[103: 96], o82_13[103: 96] };
		i82_21 <= { o82_10[ 95: 88], o82_11[ 95: 88], o82_12[ 95: 88], o82_13[ 95: 88], o82_10[ 87: 80], o82_11[ 87: 80], o82_12[ 87: 80], o82_13[ 87: 80], o82_10[ 79: 72], o82_11[ 79: 72], o82_12[ 79: 72], o82_13[ 79: 72],	o82_10[ 71: 64], o82_11[ 71: 64], o82_12[ 71: 64], o82_13[ 71: 64] };
		i82_22 <= { o82_10[ 63: 56], o82_11[ 63: 56], o82_12[ 63: 56], o82_13[ 63: 56], o82_10[ 55: 48], o82_11[ 55: 48], o82_12[ 55: 48], o82_13[ 55: 48], o82_10[ 47: 40], o82_11[ 47: 40], o82_12[ 47: 40], o82_13[ 47: 40], o82_10[ 39: 32], o82_11[ 39: 32], o82_12[ 39: 32], o82_13[ 39: 32] };
		i82_23 <= { o82_10[ 31: 24], o82_11[ 31: 24], o82_12[ 31: 24], o82_13[ 31: 24], o82_10[ 23: 16], o82_11[ 23: 16], o82_12[ 23: 16], o82_13[ 23: 16], o82_10[ 15:  8], o82_11[ 15:  8], o82_12[ 15:  8], o82_13[ 15:  8], o82_10[  7:  0], o82_11[  7:  0], o82_12[  7:  0], o82_13[  7:  0] };

	end

	reg  [127:0] i83_00, i83_01, i83_02, i83_03, i83_10, i83_11, i83_12, i83_13, i83_20, i83_21, i83_22, i83_23;
	wire [127:0] o83_00, o83_01, o83_02, o83_03, o83_10, o83_11, o83_12, o83_13, o83_20, o83_21, o83_22, o83_23;

	aes_round r83_00 (clk, i83_00, o83_00);
	aes_round r83_01 (clk, i83_01, o83_01);
	aes_round r83_02 (clk, i83_02, o83_02);
	aes_round r83_03 (clk, i83_03, o83_03);

	aes_round r83_10 (clk, i83_10, o83_10);
	aes_round r83_11 (clk, i83_11, o83_11);
	aes_round r83_12 (clk, i83_12, o83_12);
	aes_round r83_13 (clk, i83_13, o83_13);
	
	echo_mix  r83_20 (clk, i83_20, o83_20);
	echo_mix  r83_21 (clk, i83_21, o83_21);
	echo_mix  r83_22 (clk, i83_22, o83_22);
	echo_mix  r83_23 (clk, i83_23, o83_23);

	always @ ( posedge clk ) begin

		i83_00 <= { o73_20[127:120], o73_20[95:88], o73_20[63:56], o73_20[31:24], o73_21[127:120], o73_21[95:88], o73_21[63:56], o73_21[31:24], o73_22[127:120], o73_22[95:88], o73_22[63:56], o73_22[31:24], o73_23[127:120], o73_23[95:88], o73_23[63:56], o73_23[31:24] };
		i83_01 <= { o70_20[119:112], o70_20[87:80], o70_20[55:48], o70_20[23:16], o70_21[119:112], o70_21[87:80], o70_21[55:48], o70_21[23:16], o70_22[119:112], o70_22[87:80], o70_22[55:48], o70_22[23:16], o70_23[119:112], o70_23[87:80], o70_23[55:48], o70_23[23:16] };
		i83_02 <= { o71_20[111:104], o71_20[79:72], o71_20[47:40], o71_20[15: 8], o71_21[111:104], o71_21[79:72], o71_21[47:40], o71_21[15: 8], o71_22[111:104], o71_22[79:72], o71_22[47:40], o71_22[15: 8], o71_23[111:104], o71_23[79:72], o71_23[47:40], o71_23[15: 8] };
		i83_03 <= { o72_20[103: 96], o72_20[71:64], o72_20[39:32], o72_20[ 7: 0], o72_21[103: 96], o72_21[71:64], o72_21[39:32], o72_21[ 7: 0], o72_22[103: 96], o72_22[71:64], o72_22[39:32], o72_22[ 7: 0], o72_23[103: 96], o72_23[71:64], o72_23[39:32], o72_23[ 7: 0] }; 

		i83_10 <= { o83_00[127:108], o83_00[107:96] ^ 12'h028C, o83_00[95:0] };
		i83_11 <= { o83_01[127:108], o83_01[107:96] ^ 12'h0281, o83_01[95:0] };
		i83_12 <= { o83_02[127:108], o83_02[107:96] ^ 12'h0286, o83_02[95:0] };
		i83_13 <= { o83_03[127:108], o83_03[107:96] ^ 12'h028B, o83_03[95:0] };

		i83_20 <= { o83_10[127:120], o83_11[127:120], o83_12[127:120], o83_13[127:120], o83_10[119:112], o83_11[119:112], o83_12[119:112], o83_13[119:112], o83_10[111:104], o83_11[111:104], o83_12[111:104], o83_13[111:104], o83_10[103: 96], o83_11[103: 96], o83_12[103: 96], o83_13[103: 96] };
		i83_21 <= { o83_10[ 95: 88], o83_11[ 95: 88], o83_12[ 95: 88], o83_13[ 95: 88], o83_10[ 87: 80], o83_11[ 87: 80], o83_12[ 87: 80], o83_13[ 87: 80], o83_10[ 79: 72], o83_11[ 79: 72], o83_12[ 79: 72], o83_13[ 79: 72],	o83_10[ 71: 64], o83_11[ 71: 64], o83_12[ 71: 64], o83_13[ 71: 64] };
		i83_22 <= { o83_10[ 63: 56], o83_11[ 63: 56], o83_12[ 63: 56], o83_13[ 63: 56], o83_10[ 55: 48], o83_11[ 55: 48], o83_12[ 55: 48], o83_13[ 55: 48], o83_10[ 47: 40], o83_11[ 47: 40], o83_12[ 47: 40], o83_13[ 47: 40], o83_10[ 39: 32], o83_11[ 39: 32], o83_12[ 39: 32], o83_13[ 39: 32] };
		i83_23 <= { o83_10[ 31: 24], o83_11[ 31: 24], o83_12[ 31: 24], o83_13[ 31: 24], o83_10[ 23: 16], o83_11[ 23: 16], o83_12[ 23: 16], o83_13[ 23: 16], o83_10[ 15:  8], o83_11[ 15:  8], o83_12[ 15:  8], o83_13[ 15:  8], o83_10[  7:  0], o83_11[  7:  0], o83_12[  7:  0], o83_13[  7:  0] };

	end

	// ROUND 9

	reg  [127:0] i90_00, i90_01, i90_02, i90_03, i90_10, i90_11, i90_12, i90_13, i90_20, i90_21, i90_22, i90_23;
	wire [127:0] o90_00, o90_01, o90_02, o90_03, o90_10, o90_11, o90_12, o90_13, o90_20, o90_21, o90_22, o90_23;

	aes_round r90_00 (clk, i90_00, o90_00);
	aes_round r90_01 (clk, i90_01, o90_01);
	aes_round r90_02 (clk, i90_02, o90_02);
	aes_round r90_03 (clk, i90_03, o90_03);

	aes_round r90_10 (clk, i90_10, o90_10);
	aes_round r90_11 (clk, i90_11, o90_11);
	aes_round r90_12 (clk, i90_12, o90_12);
	aes_round r90_13 (clk, i90_13, o90_13);
	
	echo_mix  r90_20 (clk, i90_20, o90_20);
	echo_mix  r90_21 (clk, i90_21, o90_21);
	echo_mix  r90_22 (clk, i90_22, o90_22);
	echo_mix  r90_23 (clk, i90_23, o90_23);

	always @ ( posedge clk ) begin

		i90_00 <= { o80_20[127:120], o80_20[95:88], o80_20[63:56], o80_20[31:24], o80_21[127:120], o80_21[95:88], o80_21[63:56], o80_21[31:24], o80_22[127:120], o80_22[95:88], o80_22[63:56], o80_22[31:24], o80_23[127:120], o80_23[95:88], o80_23[63:56], o80_23[31:24] };
		i90_01 <= { o81_20[119:112], o81_20[87:80], o81_20[55:48], o81_20[23:16], o81_21[119:112], o81_21[87:80], o81_21[55:48], o81_21[23:16], o81_22[119:112], o81_22[87:80], o81_22[55:48], o81_22[23:16], o81_23[119:112], o81_23[87:80], o81_23[55:48], o81_23[23:16] };
		i90_02 <= { o82_20[111:104], o82_20[79:72], o82_20[47:40], o82_20[15: 8], o82_21[111:104], o82_21[79:72], o82_21[47:40], o82_21[15: 8], o82_22[111:104], o82_22[79:72], o82_22[47:40], o82_22[15: 8], o82_23[111:104], o82_23[79:72], o82_23[47:40], o82_23[15: 8] };
		i90_03 <= { o83_20[103: 96], o83_20[71:64], o83_20[39:32], o83_20[ 7: 0], o83_21[103: 96], o83_21[71:64], o83_21[39:32], o83_21[ 7: 0], o83_22[103: 96], o83_22[71:64], o83_22[39:32], o83_22[ 7: 0], o83_23[103: 96], o83_23[71:64], o83_23[39:32], o83_23[ 7: 0] }; 

		i90_10 <= { o90_00[127:108], o90_00[107:96] ^ 12'h0290, o90_00[95:0] };
		i90_11 <= { o90_01[127:108], o90_01[107:96] ^ 12'h0295, o90_01[95:0] };
		i90_12 <= { o90_02[127:108], o90_02[107:96] ^ 12'h029A, o90_02[95:0] };
		i90_13 <= { o90_03[127:108], o90_03[107:96] ^ 12'h029F, o90_03[95:0] };

		i90_20 <= { o90_10[127:120], o90_11[127:120], o90_12[127:120], o90_13[127:120], o90_10[119:112], o90_11[119:112], o90_12[119:112], o90_13[119:112], o90_10[111:104], o90_11[111:104], o90_12[111:104], o90_13[111:104], o90_10[103: 96], o90_11[103: 96], o90_12[103: 96], o90_13[103: 96] };
		i90_21 <= { o90_10[ 95: 88], o90_11[ 95: 88], o90_12[ 95: 88], o90_13[ 95: 88], o90_10[ 87: 80], o90_11[ 87: 80], o90_12[ 87: 80], o90_13[ 87: 80], o90_10[ 79: 72], o90_11[ 79: 72], o90_12[ 79: 72], o90_13[ 79: 72],	o90_10[ 71: 64], o90_11[ 71: 64], o90_12[ 71: 64], o90_13[ 71: 64] };
		i90_22 <= { o90_10[ 63: 56], o90_11[ 63: 56], o90_12[ 63: 56], o90_13[ 63: 56], o90_10[ 55: 48], o90_11[ 55: 48], o90_12[ 55: 48], o90_13[ 55: 48], o90_10[ 47: 40], o90_11[ 47: 40], o90_12[ 47: 40], o90_13[ 47: 40], o90_10[ 39: 32], o90_11[ 39: 32], o90_12[ 39: 32], o90_13[ 39: 32] };
		i90_23 <= { o90_10[ 31: 24], o90_11[ 31: 24], o90_12[ 31: 24], o90_13[ 31: 24], o90_10[ 23: 16], o90_11[ 23: 16], o90_12[ 23: 16], o90_13[ 23: 16], o90_10[ 15:  8], o90_11[ 15:  8], o90_12[ 15:  8], o90_13[ 15:  8], o90_10[  7:  0], o90_11[  7:  0], o90_12[  7:  0], o90_13[  7:  0] };
		
	end

//	reg  [127:0] i91_00, i91_01, i91_02, i91_03, i91_10, i91_11, i91_12, i91_13, i91_20, i91_21, i91_22, i91_23;
//	wire [127:0] o91_00, o91_01, o91_02, o91_03, o91_10, o91_11, o91_12, o91_13, o91_20, o91_21, o91_22, o91_23;
//
//	aes_round r91_00 (clk, i91_00, o91_00);
//	aes_round r91_01 (clk, i91_01, o91_01);
//	aes_round r91_02 (clk, i91_02, o91_02);
//	aes_round r91_03 (clk, i91_03, o91_03);
//
//	aes_round r91_10 (clk, i91_10, o91_10);
//	aes_round r91_11 (clk, i91_11, o91_11);
//	aes_round r91_12 (clk, i91_12, o91_12);
//	aes_round r91_13 (clk, i91_13, o91_13);
//	
//	echo_mix  r91_20 (clk, i91_20, o91_20);
//	echo_mix  r91_21 (clk, i91_21, o91_21);
//	echo_mix  r91_22 (clk, i91_22, o91_22);
//	echo_mix  r91_23 (clk, i91_23, o91_23);
//
//	always @ ( posedge clk ) begin
//
//		i91_00 <= { o81_20[127:120], o81_20[95:88], o81_20[63:56], o81_20[31:24], o81_21[127:120], o81_21[95:88], o81_21[63:56], o81_21[31:24], o81_22[127:120], o81_22[95:88], o81_22[63:56], o81_22[31:24], o81_23[127:120], o81_23[95:88], o81_23[63:56], o81_23[31:24] };
//		i91_01 <= { o82_20[119:112], o82_20[87:80], o82_20[55:48], o82_20[23:16], o82_21[119:112], o82_21[87:80], o82_21[55:48], o82_21[23:16], o82_22[119:112], o82_22[87:80], o82_22[55:48], o82_22[23:16], o82_23[119:112], o82_23[87:80], o82_23[55:48], o82_23[23:16] };
//		i91_02 <= { o83_20[111:104], o83_20[79:72], o83_20[47:40], o83_20[15: 8], o83_21[111:104], o83_21[79:72], o83_21[47:40], o83_21[15: 8], o83_22[111:104], o83_22[79:72], o83_22[47:40], o83_22[15: 8], o83_23[111:104], o83_23[79:72], o83_23[47:40], o83_23[15: 8] };
//		i91_03 <= { o80_20[103: 96], o80_20[71:64], o80_20[39:32], o80_20[ 7: 0], o80_21[103: 96], o80_21[71:64], o80_21[39:32], o80_21[ 7: 0], o80_22[103: 96], o80_22[71:64], o80_22[39:32], o80_22[ 7: 0], o80_23[103: 96], o80_23[71:64], o80_23[39:32], o80_23[ 7: 0] };
//
//		i91_10 <= { o91_00[127:108], o91_00[107:96] ^ 12'h0294, o91_00[95:0] };
//		i91_11 <= { o91_01[127:108], o91_01[107:96] ^ 12'h0299, o91_01[95:0] };
//		i91_12 <= { o91_02[127:108], o91_02[107:96] ^ 12'h029E, o91_02[95:0] };
//		i91_13 <= { o91_03[127:108], o91_03[107:96] ^ 12'h0293, o91_03[95:0] };
//
//		i91_20 <= { o91_10[127:120], o91_11[127:120], o91_12[127:120], o91_13[127:120], o91_10[119:112], o91_11[119:112], o91_12[119:112], o91_13[119:112], o91_10[111:104], o91_11[111:104], o91_12[111:104], o91_13[111:104], o91_10[103: 96], o91_11[103: 96], o91_12[103: 96], o91_13[103: 96] };
//		i91_21 <= { o91_10[ 95: 88], o91_11[ 95: 88], o91_12[ 95: 88], o91_13[ 95: 88], o91_10[ 87: 80], o91_11[ 87: 80], o91_12[ 87: 80], o91_13[ 87: 80], o91_10[ 79: 72], o91_11[ 79: 72], o91_12[ 79: 72], o91_13[ 79: 72],	o91_10[ 71: 64], o91_11[ 71: 64], o91_12[ 71: 64], o91_13[ 71: 64] };
//		i91_22 <= { o91_10[ 63: 56], o91_11[ 63: 56], o91_12[ 63: 56], o91_13[ 63: 56], o91_10[ 55: 48], o91_11[ 55: 48], o91_12[ 55: 48], o91_13[ 55: 48], o91_10[ 47: 40], o91_11[ 47: 40], o91_12[ 47: 40], o91_13[ 47: 40], o91_10[ 39: 32], o91_11[ 39: 32], o91_12[ 39: 32], o91_13[ 39: 32] };
//		i91_23 <= { o91_10[ 31: 24], o91_11[ 31: 24], o91_12[ 31: 24], o91_13[ 31: 24], o91_10[ 23: 16], o91_11[ 23: 16], o91_12[ 23: 16], o91_13[ 23: 16], o91_10[ 15:  8], o91_11[ 15:  8], o91_12[ 15:  8], o91_13[ 15:  8], o91_10[  7:  0], o91_11[  7:  0], o91_12[  7:  0], o91_13[  7:  0] };
//
//	end

	reg  [127:0] i92_00, i92_01, i92_02, i92_03, i92_10, i92_11, i92_12, i92_13, i92_20, i92_21, i92_22, i92_23;
	wire [127:0] o92_00, o92_01, o92_02, o92_03, o92_10, o92_11, o92_12, o92_13, o92_20, o92_21, o92_22, o92_23;

	aes_round r92_00 (clk, i92_00, o92_00);
	aes_round r92_01 (clk, i92_01, o92_01);
	aes_round r92_02 (clk, i92_02, o92_02);
	aes_round r92_03 (clk, i92_03, o92_03);

	aes_round r92_10 (clk, i92_10, o92_10);
	aes_round r92_11 (clk, i92_11, o92_11);
	aes_round r92_12 (clk, i92_12, o92_12);
	aes_round r92_13 (clk, i92_13, o92_13);
	
	echo_mix  r92_20 (clk, i92_20, o92_20);
	echo_mix  r92_21 (clk, i92_21, o92_21);
	echo_mix  r92_22 (clk, i92_22, o92_22);
	echo_mix  r92_23 (clk, i92_23, o92_23);

	always @ ( posedge clk ) begin

		i92_00 <= { o82_20[127:120], o82_20[95:88], o82_20[63:56], o82_20[31:24], o82_21[127:120], o82_21[95:88], o82_21[63:56], o82_21[31:24], o82_22[127:120], o82_22[95:88], o82_22[63:56], o82_22[31:24], o82_23[127:120], o82_23[95:88], o82_23[63:56], o82_23[31:24] };
		i92_01 <= { o83_20[119:112], o83_20[87:80], o83_20[55:48], o83_20[23:16], o83_21[119:112], o83_21[87:80], o83_21[55:48], o83_21[23:16], o83_22[119:112], o83_22[87:80], o83_22[55:48], o83_22[23:16], o83_23[119:112], o83_23[87:80], o83_23[55:48], o83_23[23:16] };
		i92_02 <= { o80_20[111:104], o80_20[79:72], o80_20[47:40], o80_20[15: 8], o80_21[111:104], o80_21[79:72], o80_21[47:40], o80_21[15: 8], o80_22[111:104], o80_22[79:72], o80_22[47:40], o80_22[15: 8], o80_23[111:104], o80_23[79:72], o80_23[47:40], o80_23[15: 8] };
		i92_03 <= { o81_20[103: 96], o81_20[71:64], o81_20[39:32], o81_20[ 7: 0], o81_21[103: 96], o81_21[71:64], o81_21[39:32], o81_21[ 7: 0], o81_22[103: 96], o81_22[71:64], o81_22[39:32], o81_22[ 7: 0], o81_23[103: 96], o81_23[71:64], o81_23[39:32], o81_23[ 7: 0] }; 

		i92_10 <= { o92_00[127:108], o92_00[107:96] ^ 12'h0298, o92_00[95:0] };
		i92_11 <= { o92_01[127:108], o92_01[107:96] ^ 12'h029D, o92_01[95:0] };
		i92_12 <= { o92_02[127:108], o92_02[107:96] ^ 12'h0292, o92_02[95:0] };
		i92_13 <= { o92_03[127:108], o92_03[107:96] ^ 12'h0297, o92_03[95:0] };

		i92_20 <= { o92_10[127:120], o92_11[127:120], o92_12[127:120], o92_13[127:120], o92_10[119:112], o92_11[119:112], o92_12[119:112], o92_13[119:112], o92_10[111:104], o92_11[111:104], o92_12[111:104], o92_13[111:104], o92_10[103: 96], o92_11[103: 96], o92_12[103: 96], o92_13[103: 96] };
		i92_21 <= { o92_10[ 95: 88], o92_11[ 95: 88], o92_12[ 95: 88], o92_13[ 95: 88], o92_10[ 87: 80], o92_11[ 87: 80], o92_12[ 87: 80], o92_13[ 87: 80], o92_10[ 79: 72], o92_11[ 79: 72], o92_12[ 79: 72], o92_13[ 79: 72],	o92_10[ 71: 64], o92_11[ 71: 64], o92_12[ 71: 64], o92_13[ 71: 64] };
		i92_22 <= { o92_10[ 63: 56], o92_11[ 63: 56], o92_12[ 63: 56], o92_13[ 63: 56], o92_10[ 55: 48], o92_11[ 55: 48], o92_12[ 55: 48], o92_13[ 55: 48], o92_10[ 47: 40], o92_11[ 47: 40], o92_12[ 47: 40], o92_13[ 47: 40], o92_10[ 39: 32], o92_11[ 39: 32], o92_12[ 39: 32], o92_13[ 39: 32] };
		i92_23 <= { o92_10[ 31: 24], o92_11[ 31: 24], o92_12[ 31: 24], o92_13[ 31: 24], o92_10[ 23: 16], o92_11[ 23: 16], o92_12[ 23: 16], o92_13[ 23: 16], o92_10[ 15:  8], o92_11[ 15:  8], o92_12[ 15:  8], o92_13[ 15:  8], o92_10[  7:  0], o92_11[  7:  0], o92_12[  7:  0], o92_13[  7:  0] };

	end

//	reg  [127:0] i93_00, i93_01, i93_02, i93_03, i93_10, i93_11, i93_12, i93_13, i93_20, i93_21, i93_22, i93_23;
//	wire [127:0] o93_00, o93_01, o93_02, o93_03, o93_10, o93_11, o93_12, o93_13, o93_20, o93_21, o93_22, o93_23;
//
//	aes_round r93_00 (clk, i93_00, o93_00);
//	aes_round r93_01 (clk, i93_01, o93_01);
//	aes_round r93_02 (clk, i93_02, o93_02);
//	aes_round r93_03 (clk, i93_03, o93_03);
//
//	aes_round r93_10 (clk, i93_10, o93_10);
//	aes_round r93_11 (clk, i93_11, o93_11);
//	aes_round r93_12 (clk, i93_12, o93_12);
//	aes_round r93_13 (clk, i93_13, o93_13);
//	
//	echo_mix  r93_20 (clk, i93_20, o93_20);
//	echo_mix  r93_21 (clk, i93_21, o93_21);
//	echo_mix  r93_22 (clk, i93_22, o93_22);
//	echo_mix  r93_23 (clk, i93_23, o93_23);
//
//	always @ ( posedge clk ) begin
//
//		i93_00 <= { o83_20[127:120], o83_20[95:88], o83_20[63:56], o83_20[31:24], o83_21[127:120], o83_21[95:88], o83_21[63:56], o83_21[31:24], o83_22[127:120], o83_22[95:88], o83_22[63:56], o83_22[31:24], o83_23[127:120], o83_23[95:88], o83_23[63:56], o83_23[31:24] };
//		i93_01 <= { o80_20[119:112], o80_20[87:80], o80_20[55:48], o80_20[23:16], o80_21[119:112], o80_21[87:80], o80_21[55:48], o80_21[23:16], o80_22[119:112], o80_22[87:80], o80_22[55:48], o80_22[23:16], o80_23[119:112], o80_23[87:80], o80_23[55:48], o80_23[23:16] };
//		i93_02 <= { o81_20[111:104], o81_20[79:72], o81_20[47:40], o81_20[15: 8], o81_21[111:104], o81_21[79:72], o81_21[47:40], o81_21[15: 8], o81_22[111:104], o81_22[79:72], o81_22[47:40], o81_22[15: 8], o81_23[111:104], o81_23[79:72], o81_23[47:40], o81_23[15: 8] };
//		i93_03 <= { o82_20[103: 96], o82_20[71:64], o82_20[39:32], o82_20[ 7: 0], o82_21[103: 96], o82_21[71:64], o82_21[39:32], o82_21[ 7: 0], o82_22[103: 96], o82_22[71:64], o82_22[39:32], o82_22[ 7: 0], o82_23[103: 96], o82_23[71:64], o82_23[39:32], o82_23[ 7: 0] }; 
//
//		i93_10 <= { o93_00[127:108], o93_00[107:96] ^ 12'h029C, o93_00[95:0] };
//		i93_11 <= { o93_01[127:108], o93_01[107:96] ^ 12'h0291, o93_01[95:0] };
//		i93_12 <= { o93_02[127:108], o93_02[107:96] ^ 12'h0296, o93_02[95:0] };
//		i93_13 <= { o93_03[127:108], o93_03[107:96] ^ 12'h029B, o93_03[95:0] };
//
//		i93_20 <= { o93_10[127:120], o93_11[127:120], o93_12[127:120], o93_13[127:120], o93_10[119:112], o93_11[119:112], o93_12[119:112], o93_13[119:112], o93_10[111:104], o93_11[111:104], o93_12[111:104], o93_13[111:104], o93_10[103: 96], o93_11[103: 96], o93_12[103: 96], o93_13[103: 96] };
//		i93_21 <= { o93_10[ 95: 88], o93_11[ 95: 88], o93_12[ 95: 88], o93_13[ 95: 88], o93_10[ 87: 80], o93_11[ 87: 80], o93_12[ 87: 80], o93_13[ 87: 80], o93_10[ 79: 72], o93_11[ 79: 72], o93_12[ 79: 72], o93_13[ 79: 72],	o93_10[ 71: 64], o93_11[ 71: 64], o93_12[ 71: 64], o93_13[ 71: 64] };
//		i93_22 <= { o93_10[ 63: 56], o93_11[ 63: 56], o93_12[ 63: 56], o93_13[ 63: 56], o93_10[ 55: 48], o93_11[ 55: 48], o93_12[ 55: 48], o93_13[ 55: 48], o93_10[ 47: 40], o93_11[ 47: 40], o93_12[ 47: 40], o93_13[ 47: 40], o93_10[ 39: 32], o93_11[ 39: 32], o93_12[ 39: 32], o93_13[ 39: 32] };
//		i93_23 <= { o93_10[ 31: 24], o93_11[ 31: 24], o93_12[ 31: 24], o93_13[ 31: 24], o93_10[ 23: 16], o93_11[ 23: 16], o93_12[ 23: 16], o93_13[ 23: 16], o93_10[ 15:  8], o93_11[ 15:  8], o93_12[ 15:  8], o93_13[ 15:  8], o93_10[  7:  0], o93_11[  7:  0], o93_12[  7:  0], o93_13[  7:  0] };
//
//	end


	reg [31:0] m00,m01,m02,m03,m04,m05,m06,m07,m08,m09;
	reg [31:0] m10,m11,m12,m13,m14,m15,m16,m17,m18,m19;
	reg [31:0] m20,m21,m22,m23,m24,m25,m26,m27,m28,m29;
	reg [31:0] m30,m31,m32,m33,m34,m35,m36,m37,m38,m39;
	reg [31:0] m40,m41,m42,m43,m44,m45,m46,m47,m48,m49;
	reg [31:0] m50,m51,m52,m53,m54,m55,m56,m57,m58,m59;
	reg [31:0] m60,m61,m62,m63,m64,m65,m66,m67,m68,m69;
	reg [31:0] m70,m71,m72,m73,m74,m75,m76,m77,m78,m79;
	reg [31:0] m80,m81,m82,m83,m84,m85,m86,m87,m88,m89;
	reg [31:0] m90,m91,m92,m93,m94,m95,m96,m97,m98,m99;
	reg [31:0] mA0,mA1,mA2,mA3,mA4,mA5,mA6,mA7,mA8,mA9;
	reg [31:0] mB0,mB1,mB2,mB3,mB4,mB5,mB6,mB7,mB8,mB9;
	reg [31:0] mC0,mC1,mC2,mC3,mC4,mC5,mC6,mC7,mC8,mC9;
	reg [31:0] mD0,mD1,mD2,mD3,mD4,mD5,mD6,mD7,mD8,mD9;
	reg [31:0] mE0,mE1,mE2,mE3,mE4,mE5,mE6,mE7,mE8,mE9;
	reg [31:0] mF0,mF1,mF2,mF3,mF4,mF5,mF6,mF7,mF8,mF9;

//	reg [127:0] A0_00, A0_01, A0_02, A0_03;
//	reg [127:0] A2_00, A2_01, A2_02, A2_03;

	reg [31:0] A0, A2;
	
	always @ ( posedge clk ) begin

//		A0_00 <= { o90_20[103: 96], o90_20[71:64], o90_20[39:32], o90_20[ 7: 0], o90_21[103: 96], o90_21[71:64], o90_21[39:32], o90_21[ 7: 0], o90_22[103: 96], o90_22[71:64], o90_22[39:32], o90_22[ 7: 0], o90_23[103: 96], o90_23[71:64], o90_23[39:32], o90_23[ 7: 0] };
//		A0_01 <= { o90_20[111:104], o90_20[79:72], o90_20[47:40], o90_20[15: 8], o90_21[111:104], o90_21[79:72], o90_21[47:40], o90_21[15: 8], o90_22[111:104], o90_22[79:72], o90_22[47:40], o90_22[15: 8], o90_23[111:104], o90_23[79:72], o90_23[47:40], o90_23[15: 8] };
//		A0_02 <= { o90_20[119:112], o90_20[87:80], o90_20[55:48], o90_20[23:16], o90_21[119:112], o90_21[87:80], o90_21[55:48], o90_21[23:16], o90_22[119:112], o90_22[87:80], o90_22[55:48], o90_22[23:16], o90_23[119:112], o90_23[87:80], o90_23[55:48], o90_23[23:16] }; 
//		A0_03 <= { o90_20[127:120], o90_20[95:88], o90_20[63:56], o90_20[31:24], o90_21[127:120], o90_21[95:88], o90_21[63:56], o90_21[31:24], o90_22[127:120], o90_22[95:88], o90_22[63:56], o90_22[31:24], o90_23[127:120], o90_23[95:88], o90_23[63:56], o90_23[31:24] };
//
//		A2_00 <= { o92_20[103: 96], o92_20[71:64], o92_20[39:32], o92_20[ 7: 0], o92_21[103: 96], o92_21[71:64], o92_21[39:32], o92_21[ 7: 0], o92_22[103: 96], o92_22[71:64], o92_22[39:32], o92_22[ 7: 0], o92_23[103: 96], o92_23[71:64], o92_23[39:32], o92_23[ 7: 0] };
//		A2_01 <= { o92_20[111:104], o92_20[79:72], o92_20[47:40], o92_20[15: 8], o92_21[111:104], o92_21[79:72], o92_21[47:40], o92_21[15: 8], o92_22[111:104], o92_22[79:72], o92_22[47:40], o92_22[15: 8], o92_23[111:104], o92_23[79:72], o92_23[47:40], o92_23[15: 8] };
//		A2_02 <= { o92_20[119:112], o92_20[87:80], o92_20[55:48], o92_20[23:16], o92_21[119:112], o92_21[87:80], o92_21[55:48], o92_21[23:16], o92_22[119:112], o92_22[87:80], o92_22[55:48], o92_22[23:16], o92_23[119:112], o92_23[87:80], o92_23[55:48], o92_23[23:16] }; 
//		A2_03 <= { o92_20[127:120], o92_20[95:88], o92_20[63:56], o92_20[31:24], o92_21[127:120], o92_21[95:88], o92_21[63:56], o92_21[31:24], o92_22[127:120], o92_22[95:88], o92_22[63:56], o92_22[31:24], o92_23[127:120], o92_23[95:88], o92_23[63:56], o92_23[31:24] };

		A0 <= { o90_23[119:112], o90_23[87:80], o90_23[55:48], o90_23[23:16] }; 
		A2 <= { o92_23[119:112], o92_23[87:80], o92_23[55:48], o92_23[23:16] }; 
		
		h <= A0 ^ A2 ^ mD0;

		mD9 <= mD8;
		mD8 <= mD7;
		mD7 <= mD6;
		mD6 <= mD5;
		mD5 <= mD4;
		mD4 <= mD3;
		mD3 <= mD2;
		mD2 <= mD1;
		mD1 <= mD0;
		mD0 <= mC9;
		mC9 <= mC8;
		mC8 <= mC7;
		mC7 <= mC6;
		mC6 <= mC5;
		mC5 <= mC4;
		mC4 <= mC3;
		mC3 <= mC2;
		mC2 <= mC1;
		mC1 <= mC0;
		mC0 <= mB9;
		mB9 <= mB8;
		mB8 <= mB7;
		mB7 <= mB6;
		mB6 <= mB5;
		mB5 <= mB4;
		mB4 <= mB3;
		mB3 <= mB2;
		mB2 <= mB1;
		mB1 <= mB0;
		mB0 <= mA9;
		mA9 <= mA8;
		mA8 <= mA7;
		mA7 <= mA6;
		mA6 <= mA5;
		mA5 <= mA4;
		mA4 <= mA3;
		mA3 <= mA2;
		mA2 <= mA1;
		mA1 <= mA0;
		mA0 <= m99;
		m99 <= m98;
		m98 <= m97;
		m97 <= m96;
		m96 <= m95;
		m95 <= m94;
		m94 <= m93;
		m93 <= m92;
		m92 <= m91;
		m91 <= m90;
		m90 <= m89;
		m89 <= m88;
		m88 <= m87;
		m87 <= m86;
		m86 <= m85;
		m85 <= m84;
		m84 <= m83;
		m83 <= m82;
		m82 <= m81;
		m81 <= m80;
		m80 <= m79;
		m79 <= m78;
		m78 <= m77;
		m77 <= m76;
		m76 <= m75;
		m75 <= m74;
		m74 <= m73;
		m73 <= m72;
		m72 <= m71;
		m71 <= m70;
		m70 <= m69;
		m69 <= m68;
		m68 <= m67;
		m67 <= m66;
		m66 <= m65;
		m65 <= m64;
		m64 <= m63;
		m63 <= m62;
		m62 <= m61;
		m61 <= m60;
		m60 <= m59;
		m59 <= m58;
		m58 <= m57;
		m57 <= m56;
		m56 <= m55;
		m55 <= m54;
		m54 <= m53;
		m53 <= m52;
		m52 <= m51;
		m51 <= m50;
		m50 <= m49;
		m49 <= m48;
		m48 <= m47;
		m47 <= m46;
		m46 <= m45;
		m45 <= m44;
		m44 <= m43;
		m43 <= m42;
		m42 <= m41;
		m41 <= m40;
		m40 <= m39;
		m39 <= m38;
		m38 <= m37;
		m37 <= m36;
		m36 <= m35;
		m35 <= m34;
		m34 <= m33;
		m33 <= m32;
		m32 <= m31;
		m31 <= m30;
		m30 <= m29;
		m29 <= m28;
		m28 <= m27;
		m27 <= m26;
		m26 <= m25;
		m25 <= m24;
		m24 <= m23;
		m23 <= m22;
		m22 <= m21;
		m21 <= m20;
		m20 <= m19;
		m19 <= m18;
		m18 <= m17;
		m17 <= m16;
		m16 <= m15;
		m15 <= m14;
		m14 <= m13;
		m13 <= m12;
		m12 <= m11;
		m11 <= m10;
		m10 <= m09;
		m09 <= m08;
		m08 <= m07;
		m07 <= m06;
		m06 <= m05;
		m05 <= m04;
		m04 <= m03;
		m03 <= m02;
		m02 <= m01;
		m01 <= m00;
		m00 <= msg[255:224];
		
		msg[  7:  0] <= data[511:504];
		msg[ 15:  8] <= data[503:496];
		msg[ 23: 16] <= data[495:488];
		msg[ 31: 24] <= data[487:480];
		msg[ 39: 32] <= data[479:472];
		msg[ 47: 40] <= data[471:464];
		msg[ 55: 48] <= data[463:456];
		msg[ 63: 56] <= data[455:448];
		msg[ 71: 64] <= data[447:440];
		msg[ 79: 72] <= data[439:432];
		msg[ 87: 80] <= data[431:424];
		msg[ 95: 88] <= data[423:416];
		msg[103: 96] <= data[415:408];
		msg[111:104] <= data[407:400];
		msg[119:112] <= data[399:392];
		msg[127:120] <= data[391:384];
		msg[135:128] <= data[383:376];
		msg[143:136] <= data[375:368];
		msg[151:144] <= data[367:360];
		msg[159:152] <= data[359:352];
		msg[167:160] <= data[351:344];
		msg[175:168] <= data[343:336];
		msg[183:176] <= data[335:328];
		msg[191:184] <= data[327:320];
		msg[199:192] <= data[319:312];
		msg[207:200] <= data[311:304];
		msg[215:208] <= data[303:296];
		msg[223:216] <= data[295:288];
		msg[231:224] <= data[287:280];
		msg[239:232] <= data[279:272];
		msg[247:240] <= data[271:264];
		msg[255:248] <= data[263:256];
		msg[263:256] <= data[255:248];
		msg[271:264] <= data[247:240];
		msg[279:272] <= data[239:232];
		msg[287:280] <= data[231:224];
		msg[295:288] <= data[223:216];
		msg[303:296] <= data[215:208];
		msg[311:304] <= data[207:200];
		msg[319:312] <= data[199:192];
		msg[327:320] <= data[191:184];
		msg[335:328] <= data[183:176];
		msg[343:336] <= data[175:168];
		msg[351:344] <= data[167:160];
		msg[359:352] <= data[159:152];
		msg[367:360] <= data[151:144];
		msg[375:368] <= data[143:136];
		msg[383:376] <= data[135:128];
		msg[391:384] <= data[127:120];
		msg[399:392] <= data[119:112];
		msg[407:400] <= data[111:104];
		msg[415:408] <= data[103: 96];
		msg[423:416] <= data[ 95: 88];
		msg[431:424] <= data[ 87: 80];
		msg[439:432] <= data[ 79: 72];
		msg[447:440] <= data[ 71: 64];
		msg[455:448] <= data[ 63: 56];
		msg[463:456] <= data[ 55: 48];
		msg[471:464] <= data[ 47: 40];
		msg[479:472] <= data[ 39: 32];
		msg[487:480] <= data[ 31: 24];
		msg[495:488] <= data[ 23: 16];
		msg[503:496] <= data[ 15:  8];
		msg[511:504] <= data[  7:  0];

	end
			
endmodule

module echo_mix (
	input clk,
	input [127:0] in,
	output reg [127:0] out
);

	reg [7:0] ax00, ax01, ax02, ax03;
	reg [7:0] ax10, ax11, ax12, ax13;
	reg [7:0] ax20, ax21, ax22, ax23;
	reg [7:0] ax30, ax31, ax32, ax33;

//	assign { ax03, ax02, ax01, ax00 } = in[127:96];
//	assign { ax13, ax12, ax11, ax10 } = in[ 95:64];
//	assign { ax23, ax22, ax21, ax20 } = in[ 63:32];
//	assign { ax33, ax32, ax31, ax30 } = in[ 31: 0];

	wire [7:0] a00, a01, a02, a03;
	wire [7:0] a10, a11, a12, a13;
	wire [7:0] a20, a21, a22, a23;
	wire [7:0] a30, a31, a32, a33;

	wire [7:0] b00, b01, b02, b03;
	wire [7:0] b10, b11, b12, b13;
	wire [7:0] b20, b21, b22, b23;
	wire [7:0] b30, b31, b32, b33;

	assign a00 = ax00;
	assign a01 = ax01;
	assign a02 = ax02;
	assign a03 = ax03;

	assign a10 = ax10;
	assign a11 = ax11;
	assign a12 = ax12;
	assign a13 = ax13;

	assign a20 = ax20;
	assign a21 = ax21;
	assign a22 = ax22;
	assign a23 = ax23;

	assign a30 = ax30;
	assign a31 = ax31;
	assign a32 = ax32;
	assign a33 = ax33;

	assign b00 = ax00 ^ ax03;
	assign b01 = ax01 ^ ax00;
	assign b02 = ax02 ^ ax01;
	assign b03 = ax03 ^ ax02;

	assign b10 = ax10 ^ ax13;
	assign b11 = ax11 ^ ax10;
	assign b12 = ax12 ^ ax11;
	assign b13 = ax13 ^ ax12;

	assign b20 = ax20 ^ ax23;
	assign b21 = ax21 ^ ax20;
	assign b22 = ax22 ^ ax21;
	assign b23 = ax23 ^ ax22;

	assign b30 = ax30 ^ ax33;
	assign b31 = ax31 ^ ax30;
	assign b32 = ax32 ^ ax31;
	assign b33 = ax33 ^ ax32;

//	reg [7:0] a00, a01, a02, a03;
//	reg [7:0] a10, a11, a12, a13;
//	reg [7:0] a20, a21, a22, a23;
//	reg [7:0] a30, a31, a32, a33;
//
//	reg [7:0] b00, b01, b02, b03;
//	reg [7:0] b10, b11, b12, b13;
//	reg [7:0] b20, b21, b22, b23;
//	reg [7:0] b30, b31, b32, b33;

	always @ ( posedge clk ) begin

	{ ax03, ax02, ax01, ax00 } <= in[127:96];
	{ ax13, ax12, ax11, ax10 } <= in[ 95:64];
	{ ax23, ax22, ax21, ax20 } <= in[ 63:32];
	{ ax33, ax32, ax31, ax30 } <= in[ 31: 0];

//		a00 <= ax00;
//		a01 <= ax01;
//		a02 <= ax02;
//		a03 <= ax03;
//
//		a10 <= ax10;
//		a11 <= ax11;
//		a12 <= ax12;
//		a13 <= ax13;
//
//		a20 <= ax20;
//		a21 <= ax21;
//		a22 <= ax22;
//		a23 <= ax23;
//
//		a30 <= ax30;
//		a31 <= ax31;
//		a32 <= ax32;
//		a33 <= ax33;
//		
//		b00 <= ax00 ^ ax03;
//		b01 <= ax01 ^ ax00;
//		b02 <= ax02 ^ ax01;
//		b03 <= ax03 ^ ax02;
//
//		b10 <= ax10 ^ ax13;
//		b11 <= ax11 ^ ax10;
//		b12 <= ax12 ^ ax11;
//		b13 <= ax13 ^ ax12;
//
//		b20 <= ax20 ^ ax23;
//		b21 <= ax21 ^ ax20;
//		b22 <= ax22 ^ ax21;
//		b23 <= ax23 ^ ax22;
//
//		b30 <= ax30 ^ ax33;
//		b31 <= ax31 ^ ax30;
//		b32 <= ax32 ^ ax31;
//		b33 <= ax33 ^ ax32;

	end
	
	reg [127:0] o;
	
	always @ ( * ) begin

		o[127:96] <= {
			a02[7] ^ b01[7] ^ b03[6],          a02[6] ^ b01[6] ^ b03[5],
			a02[5] ^ b01[5] ^ b03[4],          a02[4] ^ b01[4] ^ b03[3] ^ b03[7],
			a02[3] ^ b01[3] ^ b03[2] ^ b03[7], a02[2] ^ b01[2] ^ b03[1],
			a02[1] ^ b01[1] ^ b03[0] ^ b03[7], a02[0] ^ b01[0] ^ b03[7],
			a03[7] ^ b01[7] ^ b02[6],          a03[6] ^ b01[6] ^ b02[5],
			a03[5] ^ b01[5] ^ b02[4],          a03[4] ^ b01[4] ^ b02[3] ^ b02[7],
			a03[3] ^ b01[3] ^ b02[2] ^ b02[7], a03[2] ^ b01[2] ^ b02[1],
			a03[1] ^ b01[1] ^ b02[0] ^ b02[7], a03[0] ^ b01[0] ^ b02[7],
			a00[7] ^ b03[7] ^ b01[6],          a00[6] ^ b03[6] ^ b01[5],
			a00[5] ^ b03[5] ^ b01[4],          a00[4] ^ b03[4] ^ b01[3] ^ b01[7],
			a00[3] ^ b03[3] ^ b01[2] ^ b01[7], a00[2] ^ b03[2] ^ b01[1],
			a00[1] ^ b03[1] ^ b01[0] ^ b01[7], a00[0] ^ b03[0] ^ b01[7],
			a01[7] ^ b03[7] ^ b00[6],          a01[6] ^ b03[6] ^ b00[5],
			a01[5] ^ b03[5] ^ b00[4],          a01[4] ^ b03[4] ^ b00[3] ^ b00[7],
			a01[3] ^ b03[3] ^ b00[2] ^ b00[7], a01[2] ^ b03[2] ^ b00[1],
			a01[1] ^ b03[1] ^ b00[0] ^ b00[7], a01[0] ^ b03[0] ^ b00[7]
		};

		o[95:64] <= {
			a12[7] ^ b11[7] ^ b13[6],          a12[6] ^ b11[6] ^ b13[5],
			a12[5] ^ b11[5] ^ b13[4],          a12[4] ^ b11[4] ^ b13[3] ^ b13[7],
			a12[3] ^ b11[3] ^ b13[2] ^ b13[7], a12[2] ^ b11[2] ^ b13[1],
			a12[1] ^ b11[1] ^ b13[0] ^ b13[7], a12[0] ^ b11[0] ^ b13[7],
			a13[7] ^ b11[7] ^ b12[6],          a13[6] ^ b11[6] ^ b12[5],
			a13[5] ^ b11[5] ^ b12[4],          a13[4] ^ b11[4] ^ b12[3] ^ b12[7],
			a13[3] ^ b11[3] ^ b12[2] ^ b12[7], a13[2] ^ b11[2] ^ b12[1],
			a13[1] ^ b11[1] ^ b12[0] ^ b12[7], a13[0] ^ b11[0] ^ b12[7],
			a10[7] ^ b13[7] ^ b11[6],          a10[6] ^ b13[6] ^ b11[5],
			a10[5] ^ b13[5] ^ b11[4],          a10[4] ^ b13[4] ^ b11[3] ^ b11[7],
			a10[3] ^ b13[3] ^ b11[2] ^ b11[7], a10[2] ^ b13[2] ^ b11[1],
			a10[1] ^ b13[1] ^ b11[0] ^ b11[7], a10[0] ^ b13[0] ^ b11[7],
			a11[7] ^ b13[7] ^ b10[6],          a11[6] ^ b13[6] ^ b10[5],
			a11[5] ^ b13[5] ^ b10[4],          a11[4] ^ b13[4] ^ b10[3] ^ b10[7],
			a11[3] ^ b13[3] ^ b10[2] ^ b10[7], a11[2] ^ b13[2] ^ b10[1],
			a11[1] ^ b13[1] ^ b10[0] ^ b10[7], a11[0] ^ b13[0] ^ b10[7]
		};

		o[63:32] <= {
			a22[7] ^ b21[7] ^ b23[6],          a22[6] ^ b21[6] ^ b23[5],
			a22[5] ^ b21[5] ^ b23[4],          a22[4] ^ b21[4] ^ b23[3] ^ b23[7],
			a22[3] ^ b21[3] ^ b23[2] ^ b23[7], a22[2] ^ b21[2] ^ b23[1],
			a22[1] ^ b21[1] ^ b23[0] ^ b23[7], a22[0] ^ b21[0] ^ b23[7],
			a23[7] ^ b21[7] ^ b22[6],          a23[6] ^ b21[6] ^ b22[5],
			a23[5] ^ b21[5] ^ b22[4],          a23[4] ^ b21[4] ^ b22[3] ^ b22[7],
			a23[3] ^ b21[3] ^ b22[2] ^ b22[7], a23[2] ^ b21[2] ^ b22[1],
			a23[1] ^ b21[1] ^ b22[0] ^ b22[7], a23[0] ^ b21[0] ^ b22[7],
			a20[7] ^ b23[7] ^ b21[6],          a20[6] ^ b23[6] ^ b21[5],
			a20[5] ^ b23[5] ^ b21[4],          a20[4] ^ b23[4] ^ b21[3] ^ b21[7],
			a20[3] ^ b23[3] ^ b21[2] ^ b21[7], a20[2] ^ b23[2] ^ b21[1],
			a20[1] ^ b23[1] ^ b21[0] ^ b21[7], a20[0] ^ b23[0] ^ b21[7],
			a21[7] ^ b23[7] ^ b20[6],          a21[6] ^ b23[6] ^ b20[5],
			a21[5] ^ b23[5] ^ b20[4],          a21[4] ^ b23[4] ^ b20[3] ^ b20[7],
			a21[3] ^ b23[3] ^ b20[2] ^ b20[7], a21[2] ^ b23[2] ^ b20[1],
			a21[1] ^ b23[1] ^ b20[0] ^ b20[7], a21[0] ^ b23[0] ^ b20[7]
		};

		o[31:0] <= {
			a32[7] ^ b31[7] ^ b33[6],          a32[6] ^ b31[6] ^ b33[5],
			a32[5] ^ b31[5] ^ b33[4],          a32[4] ^ b31[4] ^ b33[3] ^ b33[7],
			a32[3] ^ b31[3] ^ b33[2] ^ b33[7], a32[2] ^ b31[2] ^ b33[1],
			a32[1] ^ b31[1] ^ b33[0] ^ b33[7], a32[0] ^ b31[0] ^ b33[7],
			a33[7] ^ b31[7] ^ b32[6],          a33[6] ^ b31[6] ^ b32[5],
			a33[5] ^ b31[5] ^ b32[4],          a33[4] ^ b31[4] ^ b32[3] ^ b32[7],
			a33[3] ^ b31[3] ^ b32[2] ^ b32[7], a33[2] ^ b31[2] ^ b32[1],
			a33[1] ^ b31[1] ^ b32[0] ^ b32[7], a33[0] ^ b31[0] ^ b32[7],
			a30[7] ^ b33[7] ^ b31[6],          a30[6] ^ b33[6] ^ b31[5],
			a30[5] ^ b33[5] ^ b31[4],          a30[4] ^ b33[4] ^ b31[3] ^ b31[7],
			a30[3] ^ b33[3] ^ b31[2] ^ b31[7], a30[2] ^ b33[2] ^ b31[1],
			a30[1] ^ b33[1] ^ b31[0] ^ b31[7], a30[0] ^ b33[0] ^ b31[7],
			a31[7] ^ b33[7] ^ b30[6],          a31[6] ^ b33[6] ^ b30[5],
			a31[5] ^ b33[5] ^ b30[4],          a31[4] ^ b33[4] ^ b30[3] ^ b30[7],
			a31[3] ^ b33[3] ^ b30[2] ^ b30[7], a31[2] ^ b33[2] ^ b30[1],
			a31[1] ^ b33[1] ^ b30[0] ^ b30[7], a31[0] ^ b33[0] ^ b30[7]
		};

	end

	always @ ( posedge clk ) begin
	
		out <= o;

	end
	
endmodule

module aes_round (
	input clk,
	input [127:0] in,
	output reg [127:0] out
);

	(* ram_style = "block" *) wire [7:0] s_box [0:255] = {
		8'h63, 8'h7C, 8'h77, 8'h7B, 8'hF2, 8'h6B, 8'h6F, 8'hC5, 8'h30, 8'h01, 8'h67, 8'h2B, 8'hFE, 8'hD7, 8'hAB, 8'h76, 
		8'hCA, 8'h82, 8'hC9, 8'h7D, 8'hFA, 8'h59, 8'h47, 8'hF0, 8'hAD, 8'hD4, 8'hA2, 8'hAF, 8'h9C, 8'hA4, 8'h72, 8'hC0, 
		8'hB7, 8'hFD, 8'h93, 8'h26, 8'h36, 8'h3F, 8'hF7, 8'hCC, 8'h34, 8'hA5, 8'hE5, 8'hF1, 8'h71, 8'hD8, 8'h31, 8'h15, 
		8'h04, 8'hC7, 8'h23, 8'hC3, 8'h18, 8'h96, 8'h05, 8'h9A, 8'h07, 8'h12, 8'h80, 8'hE2, 8'hEB, 8'h27, 8'hB2, 8'h75, 
		8'h09, 8'h83, 8'h2C, 8'h1A, 8'h1B, 8'h6E, 8'h5A, 8'hA0, 8'h52, 8'h3B, 8'hD6, 8'hB3, 8'h29, 8'hE3, 8'h2F, 8'h84, 
		8'h53, 8'hD1, 8'h00, 8'hED, 8'h20, 8'hFC, 8'hB1, 8'h5B, 8'h6A, 8'hCB, 8'hBE, 8'h39, 8'h4A, 8'h4C, 8'h58, 8'hCF, 
		8'hD0, 8'hEF, 8'hAA, 8'hFB, 8'h43, 8'h4D, 8'h33, 8'h85, 8'h45, 8'hF9, 8'h02, 8'h7F, 8'h50, 8'h3C, 8'h9F, 8'hA8, 
		8'h51, 8'hA3, 8'h40, 8'h8F, 8'h92, 8'h9D, 8'h38, 8'hF5, 8'hBC, 8'hB6, 8'hDA, 8'h21, 8'h10, 8'hFF, 8'hF3, 8'hD2, 
		8'hCD, 8'h0C, 8'h13, 8'hEC, 8'h5F, 8'h97, 8'h44, 8'h17, 8'hC4, 8'hA7, 8'h7E, 8'h3D, 8'h64, 8'h5D, 8'h19, 8'h73, 
		8'h60, 8'h81, 8'h4F, 8'hDC, 8'h22, 8'h2A, 8'h90, 8'h88, 8'h46, 8'hEE, 8'hB8, 8'h14, 8'hDE, 8'h5E, 8'h0B, 8'hDB, 
		8'hE0, 8'h32, 8'h3A, 8'h0A, 8'h49, 8'h06, 8'h24, 8'h5C, 8'hC2, 8'hD3, 8'hAC, 8'h62, 8'h91, 8'h95, 8'hE4, 8'h79, 
		8'hE7, 8'hC8, 8'h37, 8'h6D, 8'h8D, 8'hD5, 8'h4E, 8'hA9, 8'h6C, 8'h56, 8'hF4, 8'hEA, 8'h65, 8'h7A, 8'hAE, 8'h08, 
		8'hBA, 8'h78, 8'h25, 8'h2E, 8'h1C, 8'hA6, 8'hB4, 8'hC6, 8'hE8, 8'hDD, 8'h74, 8'h1F, 8'h4B, 8'hBD, 8'h8B, 8'h8A, 
		8'h70, 8'h3E, 8'hB5, 8'h66, 8'h48, 8'h03, 8'hF6, 8'h0E, 8'h61, 8'h35, 8'h57, 8'hB9, 8'h86, 8'hC1, 8'h1D, 8'h9E, 
		8'hE1, 8'hF8, 8'h98, 8'h11, 8'h69, 8'hD9, 8'h8E, 8'h94, 8'h9B, 8'h1E, 8'h87, 8'hE9, 8'hCE, 8'h55, 8'h28, 8'hDF, 
		8'h8C, 8'hA1, 8'h89, 8'h0D, 8'hBF, 8'hE6, 8'h42, 8'h68, 8'h41, 8'h99, 8'h2D, 8'h0F, 8'hB0, 8'h54, 8'hBB, 8'h16
	};

	reg [127:0] i;
			
	always @ ( posedge clk ) begin
	
		i <= in;

	end
	
	reg[7:0] sb0x,sb1x,sb2x,sb3x,sb4x,sb5x,sb6x,sb7x,sb8x,sb9x,sbAx,sbBx,sbCx,sbDx,sbEx,sbFx;
	reg[7:0] sb0,sb1,sb2,sb3,sb4,sb5,sb6,sb7,sb8,sb9,sbA,sbB,sbC,sbD,sbE,sbF;
			
	always @ ( posedge clk ) begin

		sbFx <= s_box[i[63:56]];
		sbEx <= s_box[i[95:88]];
		sbDx <= s_box[i[127:120]];
		sbCx <= s_box[i[31:24]];
		sbBx <= s_box[i[87:80]];
		sbAx <= s_box[i[119:112]];
		sb9x <= s_box[i[23:16]];
		sb8x <= s_box[i[55:48]];
		sb7x <= s_box[i[111:104]];
		sb6x <= s_box[i[15:8]];
		sb5x <= s_box[i[47:40]];
		sb4x <= s_box[i[79:72]];
		sb3x <= s_box[i[7:0]];
		sb2x <= s_box[i[39:32]];
		sb1x <= s_box[i[71:64]];
		sb0x <= s_box[i[103:96]];

		// Extra FF To Allow Use Of Block Ram Output Register
		sbF <= sbFx;
		sbE <= sbEx;
		sbD <= sbDx;
		sbC <= sbCx;
		sbB <= sbBx;
		sbA <= sbAx;
		sb9 <= sb9x;
		sb8 <= sb8x;
		sb7 <= sb7x;
		sb6 <= sb6x;
		sb5 <= sb5x;
		sb4 <= sb4x;
		sb3 <= sb3x;
		sb2 <= sb2x;
		sb1 <= sb1x;
		sb0 <= sb0x;

	end

//	reg[7:0] g1_0,g1_1,g1_2,g1_3,g1_4,g1_5,g1_6,g1_7,g1_8,g1_9,g1_A,g1_B,g1_C,g1_D,g1_E,g1_F;
//	reg[7:0] g2_0,g2_1,g2_2,g2_3,g2_4,g2_5,g2_6,g2_7,g2_8,g2_9,g2_A,g2_B,g2_C,g2_D,g2_E,g2_F;
//
//	always @ ( posedge clk ) begin
//
//		g1_0 <= sb0;
//		g1_1 <= sb1;
//		g1_2 <= sb2;
//		g1_3 <= sb3;
//		g1_4 <= sb4;
//		g1_5 <= sb5;
//		g1_6 <= sb6;
//		g1_7 <= sb7;
//		g1_8 <= sb8;
//		g1_9 <= sb9;
//		g1_A <= sbA;
//		g1_B <= sbB;
//		g1_C <= sbC;
//		g1_D <= sbD;
//		g1_E <= sbE;
//		g1_F <= sbF;
//
//		g2_0 <= gf_2(sb0);
//		g2_1 <= gf_2(sb1);
//		g2_2 <= gf_2(sb2);
//		g2_3 <= gf_2(sb3);
//		g2_4 <= gf_2(sb4);
//		g2_5 <= gf_2(sb5);
//		g2_6 <= gf_2(sb6);
//		g2_7 <= gf_2(sb7);
//		g2_8 <= gf_2(sb8);
//		g2_9 <= gf_2(sb9);
//		g2_A <= gf_2(sbA);
//		g2_B <= gf_2(sbB);
//		g2_C <= gf_2(sbC);
//		g2_D <= gf_2(sbD);
//		g2_E <= gf_2(sbE);
//		g2_F <= gf_2(sbF);
//
//	end

	wire [7:0] g1_0,g1_1,g1_2,g1_3,g1_4,g1_5,g1_6,g1_7,g1_8,g1_9,g1_A,g1_B,g1_C,g1_D,g1_E,g1_F;
	wire [7:0] g2_0,g2_1,g2_2,g2_3,g2_4,g2_5,g2_6,g2_7,g2_8,g2_9,g2_A,g2_B,g2_C,g2_D,g2_E,g2_F;
	
	assign g1_0 = sb0;
	assign g1_1 = sb1;
	assign g1_2 = sb2;
	assign g1_3 = sb3;
	assign g1_4 = sb4;
	assign g1_5 = sb5;
	assign g1_6 = sb6;
	assign g1_7 = sb7;
	assign g1_8 = sb8;
	assign g1_9 = sb9;
	assign g1_A = sbA;
	assign g1_B = sbB;
	assign g1_C = sbC;
	assign g1_D = sbD;
	assign g1_E = sbE;
	assign g1_F = sbF;

	assign g2_0 = gf_2(sb0);
	assign g2_1 = gf_2(sb1);
	assign g2_2 = gf_2(sb2);
	assign g2_3 = gf_2(sb3);
	assign g2_4 = gf_2(sb4);
	assign g2_5 = gf_2(sb5);
	assign g2_6 = gf_2(sb6);
	assign g2_7 = gf_2(sb7);
	assign g2_8 = gf_2(sb8);
	assign g2_9 = gf_2(sb9);
	assign g2_A = gf_2(sbA);
	assign g2_B = gf_2(sbB);
	assign g2_C = gf_2(sbC);
	assign g2_D = gf_2(sbD);
	assign g2_E = gf_2(sbE);
	assign g2_F = gf_2(sbF);

	reg[7:0] o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,oA,oB,oC,oD,oE,oF;

	always @ ( * ) begin
	
		o0 <= g2_C ^ g2_0 ^ g1_0 ^ g1_4 ^ g1_8;
		o1 <= g2_8 ^ g2_C ^ g1_C ^ g1_0 ^ g1_4;
		o2 <= g2_4 ^ g2_8 ^ g1_8 ^ g1_C ^ g1_0;
		o3 <= g2_0 ^ g2_4 ^ g1_4 ^ g1_8 ^ g1_C;
		o4 <= g2_D ^ g2_1 ^ g1_1 ^ g1_5 ^ g1_9;
		o5 <= g2_9 ^ g2_D ^ g1_D ^ g1_1 ^ g1_5;
		o6 <= g2_5 ^ g2_9 ^ g1_9 ^ g1_D ^ g1_1;
		o7 <= g2_1 ^ g2_5 ^ g1_5 ^ g1_9 ^ g1_D;
		o8 <= g2_E ^ g2_2 ^ g1_2 ^ g1_6 ^ g1_A;
		o9 <= g2_A ^ g2_E ^ g1_E ^ g1_2 ^ g1_6;
		oA <= g2_6 ^ g2_A ^ g1_A ^ g1_E ^ g1_2;
		oB <= g2_2 ^ g2_6 ^ g1_6 ^ g1_A ^ g1_E;
		oC <= g2_F ^ g2_3 ^ g1_3 ^ g1_7 ^ g1_B;
		oD <= g2_B ^ g2_F ^ g1_F ^ g1_3 ^ g1_7;
		oE <= g2_7 ^ g2_B ^ g1_B ^ g1_F ^ g1_3;
		oF <= g2_3 ^ g2_7 ^ g1_7 ^ g1_B ^ g1_F;
		
	end

	always @ ( posedge clk ) begin
			
		out <= { o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,oA,oB,oC,oD,oE,oF };
		
	end
			
	// Calculate GF(256) Multiplication (x2)
	function [7:0] gf_2;
		input [7:0] n;
		begin
			gf_2 = {n[6],n[5],n[4],n[3]^n[7],n[2]^n[7],n[1],n[0]^n[7],n[7]};
		end
	endfunction
	
endmodule
