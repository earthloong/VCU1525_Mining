/*
 * Copyright (c) 2016 Sprocket
 *
 * This is free software: you can redistribute it and/or modify
 * it under the terms of the GNU Affero General Public License with
 * additional permissions to the one published by the Free Software
 * Foundation, either version 3 of the License, or (at your option)
 * any later version. For more information see LICENSE.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU Affero General Public License for more details.
 *
 * You should have received a copy of the GNU Affero General Public License
 * along with this program. If not, see <http://www.gnu.org/licenses/>.
 */

module mix_bytes(
	input  clk,
	input  [1023:0] in,
	output reg [1023:0] out
);

	reg [63:0] m0, m1, m2, m3, m4, m5, m6, m7;
	reg [63:0] m8, m9, mA, mB, mC, mD, mE, mF;
	
	reg [7:0] b00,b01,b02,b03,b04,b05,b06,b07;
	reg [7:0] b00_2,b01_2,b02_2,b03_2,b04_2,b05_2,b06_2,b07_2;
	reg [7:0] b00_4,b01_4,b02_4,b03_4,b04_4,b05_4,b06_4,b07_4;

	always @ (*) begin
	
		{ b00, b01, b02, b03, b04, b05, b06, b07 } = in[1023:960];
		
		b00_2 = {b00[6], b00[5], b00[4], b00[3]^b00[7], b00[2]^b00[7], b00[1], b00[0]^b00[7], b00[7]};
		b01_2 = {b01[6], b01[5], b01[4], b01[3]^b01[7], b01[2]^b01[7], b01[1], b01[0]^b01[7], b01[7]};
		b02_2 = {b02[6], b02[5], b02[4], b02[3]^b02[7], b02[2]^b02[7], b02[1], b02[0]^b02[7], b02[7]};
		b03_2 = {b03[6], b03[5], b03[4], b03[3]^b03[7], b03[2]^b03[7], b03[1], b03[0]^b03[7], b03[7]};
		b04_2 = {b04[6], b04[5], b04[4], b04[3]^b04[7], b04[2]^b04[7], b04[1], b04[0]^b04[7], b04[7]};
		b05_2 = {b05[6], b05[5], b05[4], b05[3]^b05[7], b05[2]^b05[7], b05[1], b05[0]^b05[7], b05[7]};
		b06_2 = {b06[6], b06[5], b06[4], b06[3]^b06[7], b06[2]^b06[7], b06[1], b06[0]^b06[7], b06[7]};
		b07_2 = {b07[6], b07[5], b07[4], b07[3]^b07[7], b07[2]^b07[7], b07[1], b07[0]^b07[7], b07[7]};

		b00_4 = {b00[5], b00[4], b00[3]^ b00[7], b00[2]^ b00[7]^b00[6], b00[6]^b00[1], b00[0]^b00[7], b00[6]^b00[7], b00[6]};
		b01_4 = {b01[5], b01[4], b01[3]^ b01[7], b01[2]^ b01[7]^b01[6], b01[6]^b01[1], b01[0]^b01[7], b01[6]^b01[7], b01[6]};
		b02_4 = {b02[5], b02[4], b02[3]^ b02[7], b02[2]^ b02[7]^b02[6], b02[6]^b02[1], b02[0]^b02[7], b02[6]^b02[7], b02[6]};
		b03_4 = {b03[5], b03[4], b03[3]^ b03[7], b03[2]^ b03[7]^b03[6], b03[6]^b03[1], b03[0]^b03[7], b03[6]^b03[7], b03[6]};
		b04_4 = {b04[5], b04[4], b04[3]^ b04[7], b04[2]^ b04[7]^b04[6], b04[6]^b04[1], b04[0]^b04[7], b04[6]^b04[7], b04[6]};
		b05_4 = {b05[5], b05[4], b05[3]^ b05[7], b05[2]^ b05[7]^b05[6], b05[6]^b05[1], b05[0]^b05[7], b05[6]^b05[7], b05[6]};
		b06_4 = {b06[5], b06[4], b06[3]^ b06[7], b06[2]^ b06[7]^b06[6], b06[6]^b06[1], b06[0]^b06[7], b06[6]^b06[7], b06[6]};
		b07_4 = {b07[5], b07[4], b07[3]^ b07[7], b07[2]^ b07[7]^b07[6], b07[6]^b07[1], b07[0]^b07[7], b07[6]^b07[7], b07[6]};

		m0 = {
			b00_2 ^ b01_2 ^ b02_2 ^ b02 ^ b03_4 ^ b04_4 ^ b04 ^ b05_2 ^ b05 ^ b06_4 ^ b06 ^ b07_4 ^ b07_2 ^ b07,
			b01_2 ^ b02_2 ^ b03_2 ^ b03 ^ b04_4 ^ b05_4 ^ b05 ^ b06_2 ^ b06 ^ b07_4 ^ b07 ^ b00_4 ^ b00_2 ^ b00,
			b02_2 ^ b03_2 ^ b04_2 ^ b04 ^ b05_4 ^ b06_4 ^ b06 ^ b07_2 ^ b07 ^ b00_4 ^ b00 ^ b01_4 ^ b01_2 ^ b01,
			b03_2 ^ b04_2 ^ b05_2 ^ b05 ^ b06_4 ^ b07_4 ^ b07 ^ b00_2 ^ b00 ^ b01_4 ^ b01 ^ b02_4 ^ b02_2 ^ b02,
			b04_2 ^ b05_2 ^ b06_2 ^ b06 ^ b07_4 ^ b00_4 ^ b00 ^ b01_2 ^ b01 ^ b02_4 ^ b02 ^ b03_4 ^ b03_2 ^ b03,
			b05_2 ^ b06_2 ^ b07_2 ^ b07 ^ b00_4 ^ b01_4 ^ b01 ^ b02_2 ^ b02 ^ b03_4 ^ b03 ^ b04_4 ^ b04_2 ^ b04,
			b06_2 ^ b07_2 ^ b00_2 ^ b00 ^ b01_4 ^ b02_4 ^ b02 ^ b03_2 ^ b03 ^ b04_4 ^ b04 ^ b05_4 ^ b05_2 ^ b05,
			b07_2 ^ b00_2 ^ b01_2 ^ b01 ^ b02_4 ^ b03_4 ^ b03 ^ b04_2 ^ b04 ^ b05_4 ^ b05 ^ b06_4 ^ b06_2 ^ b06
		};

	end

	reg [7:0] b10,b11,b12,b13,b14,b15,b16,b17;
	reg [7:0] b10_2,b11_2,b12_2,b13_2,b14_2,b15_2,b16_2,b17_2;
	reg [7:0] b10_4,b11_4,b12_4,b13_4,b14_4,b15_4,b16_4,b17_4;

	always @ (*) begin
	
		{ b10, b11, b12, b13, b14, b15, b16, b17 } = in[959:896];
		
		b10_2 = {b10[6], b10[5], b10[4], b10[3]^b10[7], b10[2]^b10[7], b10[1], b10[0]^b10[7], b10[7]};
		b11_2 = {b11[6], b11[5], b11[4], b11[3]^b11[7], b11[2]^b11[7], b11[1], b11[0]^b11[7], b11[7]};
		b12_2 = {b12[6], b12[5], b12[4], b12[3]^b12[7], b12[2]^b12[7], b12[1], b12[0]^b12[7], b12[7]};
		b13_2 = {b13[6], b13[5], b13[4], b13[3]^b13[7], b13[2]^b13[7], b13[1], b13[0]^b13[7], b13[7]};
		b14_2 = {b14[6], b14[5], b14[4], b14[3]^b14[7], b14[2]^b14[7], b14[1], b14[0]^b14[7], b14[7]};
		b15_2 = {b15[6], b15[5], b15[4], b15[3]^b15[7], b15[2]^b15[7], b15[1], b15[0]^b15[7], b15[7]};
		b16_2 = {b16[6], b16[5], b16[4], b16[3]^b16[7], b16[2]^b16[7], b16[1], b16[0]^b16[7], b16[7]};
		b17_2 = {b17[6], b17[5], b17[4], b17[3]^b17[7], b17[2]^b17[7], b17[1], b17[0]^b17[7], b17[7]};

		b10_4 = {b10[5], b10[4], b10[3]^ b10[7], b10[2]^ b10[7]^b10[6], b10[6]^b10[1], b10[0]^b10[7], b10[6]^b10[7], b10[6]};
		b11_4 = {b11[5], b11[4], b11[3]^ b11[7], b11[2]^ b11[7]^b11[6], b11[6]^b11[1], b11[0]^b11[7], b11[6]^b11[7], b11[6]};
		b12_4 = {b12[5], b12[4], b12[3]^ b12[7], b12[2]^ b12[7]^b12[6], b12[6]^b12[1], b12[0]^b12[7], b12[6]^b12[7], b12[6]};
		b13_4 = {b13[5], b13[4], b13[3]^ b13[7], b13[2]^ b13[7]^b13[6], b13[6]^b13[1], b13[0]^b13[7], b13[6]^b13[7], b13[6]};
		b14_4 = {b14[5], b14[4], b14[3]^ b14[7], b14[2]^ b14[7]^b14[6], b14[6]^b14[1], b14[0]^b14[7], b14[6]^b14[7], b14[6]};
		b15_4 = {b15[5], b15[4], b15[3]^ b15[7], b15[2]^ b15[7]^b15[6], b15[6]^b15[1], b15[0]^b15[7], b15[6]^b15[7], b15[6]};
		b16_4 = {b16[5], b16[4], b16[3]^ b16[7], b16[2]^ b16[7]^b16[6], b16[6]^b16[1], b16[0]^b16[7], b16[6]^b16[7], b16[6]};
		b17_4 = {b17[5], b17[4], b17[3]^ b17[7], b17[2]^ b17[7]^b17[6], b17[6]^b17[1], b17[0]^b17[7], b17[6]^b17[7], b17[6]};

		m1 = {
			b10_2 ^ b11_2 ^ b12_2 ^ b12 ^ b13_4 ^ b14_4 ^ b14 ^ b15_2 ^ b15 ^ b16_4 ^ b16 ^ b17_4 ^ b17_2 ^ b17,
			b11_2 ^ b12_2 ^ b13_2 ^ b13 ^ b14_4 ^ b15_4 ^ b15 ^ b16_2 ^ b16 ^ b17_4 ^ b17 ^ b10_4 ^ b10_2 ^ b10,
			b12_2 ^ b13_2 ^ b14_2 ^ b14 ^ b15_4 ^ b16_4 ^ b16 ^ b17_2 ^ b17 ^ b10_4 ^ b10 ^ b11_4 ^ b11_2 ^ b11,
			b13_2 ^ b14_2 ^ b15_2 ^ b15 ^ b16_4 ^ b17_4 ^ b17 ^ b10_2 ^ b10 ^ b11_4 ^ b11 ^ b12_4 ^ b12_2 ^ b12,
			b14_2 ^ b15_2 ^ b16_2 ^ b16 ^ b17_4 ^ b10_4 ^ b10 ^ b11_2 ^ b11 ^ b12_4 ^ b12 ^ b13_4 ^ b13_2 ^ b13,
			b15_2 ^ b16_2 ^ b17_2 ^ b17 ^ b10_4 ^ b11_4 ^ b11 ^ b12_2 ^ b12 ^ b13_4 ^ b13 ^ b14_4 ^ b14_2 ^ b14,
			b16_2 ^ b17_2 ^ b10_2 ^ b10 ^ b11_4 ^ b12_4 ^ b12 ^ b13_2 ^ b13 ^ b14_4 ^ b14 ^ b15_4 ^ b15_2 ^ b15,
			b17_2 ^ b10_2 ^ b11_2 ^ b11 ^ b12_4 ^ b13_4 ^ b13 ^ b14_2 ^ b14 ^ b15_4 ^ b15 ^ b16_4 ^ b16_2 ^ b16
		};

	end

	reg [7:0] b20,b21,b22,b23,b24,b25,b26,b27;
	reg [7:0] b20_2,b21_2,b22_2,b23_2,b24_2,b25_2,b26_2,b27_2;
	reg [7:0] b20_4,b21_4,b22_4,b23_4,b24_4,b25_4,b26_4,b27_4;

	always @ (*) begin
	
		{ b20, b21, b22, b23, b24, b25, b26, b27 } = in[895:832];
		
		b20_2 = {b20[6], b20[5], b20[4], b20[3]^b20[7], b20[2]^b20[7], b20[1], b20[0]^b20[7], b20[7]};
		b21_2 = {b21[6], b21[5], b21[4], b21[3]^b21[7], b21[2]^b21[7], b21[1], b21[0]^b21[7], b21[7]};
		b22_2 = {b22[6], b22[5], b22[4], b22[3]^b22[7], b22[2]^b22[7], b22[1], b22[0]^b22[7], b22[7]};
		b23_2 = {b23[6], b23[5], b23[4], b23[3]^b23[7], b23[2]^b23[7], b23[1], b23[0]^b23[7], b23[7]};
		b24_2 = {b24[6], b24[5], b24[4], b24[3]^b24[7], b24[2]^b24[7], b24[1], b24[0]^b24[7], b24[7]};
		b25_2 = {b25[6], b25[5], b25[4], b25[3]^b25[7], b25[2]^b25[7], b25[1], b25[0]^b25[7], b25[7]};
		b26_2 = {b26[6], b26[5], b26[4], b26[3]^b26[7], b26[2]^b26[7], b26[1], b26[0]^b26[7], b26[7]};
		b27_2 = {b27[6], b27[5], b27[4], b27[3]^b27[7], b27[2]^b27[7], b27[1], b27[0]^b27[7], b27[7]};

		b20_4 = {b20[5], b20[4], b20[3]^ b20[7], b20[2]^ b20[7]^b20[6], b20[6]^b20[1], b20[0]^b20[7], b20[6]^b20[7], b20[6]};
		b21_4 = {b21[5], b21[4], b21[3]^ b21[7], b21[2]^ b21[7]^b21[6], b21[6]^b21[1], b21[0]^b21[7], b21[6]^b21[7], b21[6]};
		b22_4 = {b22[5], b22[4], b22[3]^ b22[7], b22[2]^ b22[7]^b22[6], b22[6]^b22[1], b22[0]^b22[7], b22[6]^b22[7], b22[6]};
		b23_4 = {b23[5], b23[4], b23[3]^ b23[7], b23[2]^ b23[7]^b23[6], b23[6]^b23[1], b23[0]^b23[7], b23[6]^b23[7], b23[6]};
		b24_4 = {b24[5], b24[4], b24[3]^ b24[7], b24[2]^ b24[7]^b24[6], b24[6]^b24[1], b24[0]^b24[7], b24[6]^b24[7], b24[6]};
		b25_4 = {b25[5], b25[4], b25[3]^ b25[7], b25[2]^ b25[7]^b25[6], b25[6]^b25[1], b25[0]^b25[7], b25[6]^b25[7], b25[6]};
		b26_4 = {b26[5], b26[4], b26[3]^ b26[7], b26[2]^ b26[7]^b26[6], b26[6]^b26[1], b26[0]^b26[7], b26[6]^b26[7], b26[6]};
		b27_4 = {b27[5], b27[4], b27[3]^ b27[7], b27[2]^ b27[7]^b27[6], b27[6]^b27[1], b27[0]^b27[7], b27[6]^b27[7], b27[6]};

		m2 = {
			b20_2 ^ b21_2 ^ b22_2 ^ b22 ^ b23_4 ^ b24_4 ^ b24 ^ b25_2 ^ b25 ^ b26_4 ^ b26 ^ b27_4 ^ b27_2 ^ b27,
			b21_2 ^ b22_2 ^ b23_2 ^ b23 ^ b24_4 ^ b25_4 ^ b25 ^ b26_2 ^ b26 ^ b27_4 ^ b27 ^ b20_4 ^ b20_2 ^ b20,
			b22_2 ^ b23_2 ^ b24_2 ^ b24 ^ b25_4 ^ b26_4 ^ b26 ^ b27_2 ^ b27 ^ b20_4 ^ b20 ^ b21_4 ^ b21_2 ^ b21,
			b23_2 ^ b24_2 ^ b25_2 ^ b25 ^ b26_4 ^ b27_4 ^ b27 ^ b20_2 ^ b20 ^ b21_4 ^ b21 ^ b22_4 ^ b22_2 ^ b22,
			b24_2 ^ b25_2 ^ b26_2 ^ b26 ^ b27_4 ^ b20_4 ^ b20 ^ b21_2 ^ b21 ^ b22_4 ^ b22 ^ b23_4 ^ b23_2 ^ b23,
			b25_2 ^ b26_2 ^ b27_2 ^ b27 ^ b20_4 ^ b21_4 ^ b21 ^ b22_2 ^ b22 ^ b23_4 ^ b23 ^ b24_4 ^ b24_2 ^ b24,
			b26_2 ^ b27_2 ^ b20_2 ^ b20 ^ b21_4 ^ b22_4 ^ b22 ^ b23_2 ^ b23 ^ b24_4 ^ b24 ^ b25_4 ^ b25_2 ^ b25,
			b27_2 ^ b20_2 ^ b21_2 ^ b21 ^ b22_4 ^ b23_4 ^ b23 ^ b24_2 ^ b24 ^ b25_4 ^ b25 ^ b26_4 ^ b26_2 ^ b26
		};

	end

	reg [7:0] b30,b31,b32,b33,b34,b35,b36,b37;
	reg [7:0] b30_2,b31_2,b32_2,b33_2,b34_2,b35_2,b36_2,b37_2;
	reg [7:0] b30_4,b31_4,b32_4,b33_4,b34_4,b35_4,b36_4,b37_4;

	always @ (*) begin
	
		{ b30, b31, b32, b33, b34, b35, b36, b37 } = in[831:768];
		
		b30_2 = {b30[6], b30[5], b30[4], b30[3]^b30[7], b30[2]^b30[7], b30[1], b30[0]^b30[7], b30[7]};
		b31_2 = {b31[6], b31[5], b31[4], b31[3]^b31[7], b31[2]^b31[7], b31[1], b31[0]^b31[7], b31[7]};
		b32_2 = {b32[6], b32[5], b32[4], b32[3]^b32[7], b32[2]^b32[7], b32[1], b32[0]^b32[7], b32[7]};
		b33_2 = {b33[6], b33[5], b33[4], b33[3]^b33[7], b33[2]^b33[7], b33[1], b33[0]^b33[7], b33[7]};
		b34_2 = {b34[6], b34[5], b34[4], b34[3]^b34[7], b34[2]^b34[7], b34[1], b34[0]^b34[7], b34[7]};
		b35_2 = {b35[6], b35[5], b35[4], b35[3]^b35[7], b35[2]^b35[7], b35[1], b35[0]^b35[7], b35[7]};
		b36_2 = {b36[6], b36[5], b36[4], b36[3]^b36[7], b36[2]^b36[7], b36[1], b36[0]^b36[7], b36[7]};
		b37_2 = {b37[6], b37[5], b37[4], b37[3]^b37[7], b37[2]^b37[7], b37[1], b37[0]^b37[7], b37[7]};

		b30_4 = {b30[5], b30[4], b30[3]^ b30[7], b30[2]^ b30[7]^b30[6], b30[6]^b30[1], b30[0]^b30[7], b30[6]^b30[7], b30[6]};
		b31_4 = {b31[5], b31[4], b31[3]^ b31[7], b31[2]^ b31[7]^b31[6], b31[6]^b31[1], b31[0]^b31[7], b31[6]^b31[7], b31[6]};
		b32_4 = {b32[5], b32[4], b32[3]^ b32[7], b32[2]^ b32[7]^b32[6], b32[6]^b32[1], b32[0]^b32[7], b32[6]^b32[7], b32[6]};
		b33_4 = {b33[5], b33[4], b33[3]^ b33[7], b33[2]^ b33[7]^b33[6], b33[6]^b33[1], b33[0]^b33[7], b33[6]^b33[7], b33[6]};
		b34_4 = {b34[5], b34[4], b34[3]^ b34[7], b34[2]^ b34[7]^b34[6], b34[6]^b34[1], b34[0]^b34[7], b34[6]^b34[7], b34[6]};
		b35_4 = {b35[5], b35[4], b35[3]^ b35[7], b35[2]^ b35[7]^b35[6], b35[6]^b35[1], b35[0]^b35[7], b35[6]^b35[7], b35[6]};
		b36_4 = {b36[5], b36[4], b36[3]^ b36[7], b36[2]^ b36[7]^b36[6], b36[6]^b36[1], b36[0]^b36[7], b36[6]^b36[7], b36[6]};
		b37_4 = {b37[5], b37[4], b37[3]^ b37[7], b37[2]^ b37[7]^b37[6], b37[6]^b37[1], b37[0]^b37[7], b37[6]^b37[7], b37[6]};

		m3 = {
			b30_2 ^ b31_2 ^ b32_2 ^ b32 ^ b33_4 ^ b34_4 ^ b34 ^ b35_2 ^ b35 ^ b36_4 ^ b36 ^ b37_4 ^ b37_2 ^ b37,
			b31_2 ^ b32_2 ^ b33_2 ^ b33 ^ b34_4 ^ b35_4 ^ b35 ^ b36_2 ^ b36 ^ b37_4 ^ b37 ^ b30_4 ^ b30_2 ^ b30,
			b32_2 ^ b33_2 ^ b34_2 ^ b34 ^ b35_4 ^ b36_4 ^ b36 ^ b37_2 ^ b37 ^ b30_4 ^ b30 ^ b31_4 ^ b31_2 ^ b31,
			b33_2 ^ b34_2 ^ b35_2 ^ b35 ^ b36_4 ^ b37_4 ^ b37 ^ b30_2 ^ b30 ^ b31_4 ^ b31 ^ b32_4 ^ b32_2 ^ b32,
			b34_2 ^ b35_2 ^ b36_2 ^ b36 ^ b37_4 ^ b30_4 ^ b30 ^ b31_2 ^ b31 ^ b32_4 ^ b32 ^ b33_4 ^ b33_2 ^ b33,
			b35_2 ^ b36_2 ^ b37_2 ^ b37 ^ b30_4 ^ b31_4 ^ b31 ^ b32_2 ^ b32 ^ b33_4 ^ b33 ^ b34_4 ^ b34_2 ^ b34,
			b36_2 ^ b37_2 ^ b30_2 ^ b30 ^ b31_4 ^ b32_4 ^ b32 ^ b33_2 ^ b33 ^ b34_4 ^ b34 ^ b35_4 ^ b35_2 ^ b35,
			b37_2 ^ b30_2 ^ b31_2 ^ b31 ^ b32_4 ^ b33_4 ^ b33 ^ b34_2 ^ b34 ^ b35_4 ^ b35 ^ b36_4 ^ b36_2 ^ b36
		};

	end

	reg [7:0] b40,b41,b42,b43,b44,b45,b46,b47;
	reg [7:0] b40_2,b41_2,b42_2,b43_2,b44_2,b45_2,b46_2,b47_2;
	reg [7:0] b40_4,b41_4,b42_4,b43_4,b44_4,b45_4,b46_4,b47_4;

	always @ (*) begin
	
		{ b40, b41, b42, b43, b44, b45, b46, b47 } = in[767:704];
		
		b40_2 = {b40[6], b40[5], b40[4], b40[3]^b40[7], b40[2]^b40[7], b40[1], b40[0]^b40[7], b40[7]};
		b41_2 = {b41[6], b41[5], b41[4], b41[3]^b41[7], b41[2]^b41[7], b41[1], b41[0]^b41[7], b41[7]};
		b42_2 = {b42[6], b42[5], b42[4], b42[3]^b42[7], b42[2]^b42[7], b42[1], b42[0]^b42[7], b42[7]};
		b43_2 = {b43[6], b43[5], b43[4], b43[3]^b43[7], b43[2]^b43[7], b43[1], b43[0]^b43[7], b43[7]};
		b44_2 = {b44[6], b44[5], b44[4], b44[3]^b44[7], b44[2]^b44[7], b44[1], b44[0]^b44[7], b44[7]};
		b45_2 = {b45[6], b45[5], b45[4], b45[3]^b45[7], b45[2]^b45[7], b45[1], b45[0]^b45[7], b45[7]};
		b46_2 = {b46[6], b46[5], b46[4], b46[3]^b46[7], b46[2]^b46[7], b46[1], b46[0]^b46[7], b46[7]};
		b47_2 = {b47[6], b47[5], b47[4], b47[3]^b47[7], b47[2]^b47[7], b47[1], b47[0]^b47[7], b47[7]};

		b40_4 = {b40[5], b40[4], b40[3]^ b40[7], b40[2]^ b40[7]^b40[6], b40[6]^b40[1], b40[0]^b40[7], b40[6]^b40[7], b40[6]};
		b41_4 = {b41[5], b41[4], b41[3]^ b41[7], b41[2]^ b41[7]^b41[6], b41[6]^b41[1], b41[0]^b41[7], b41[6]^b41[7], b41[6]};
		b42_4 = {b42[5], b42[4], b42[3]^ b42[7], b42[2]^ b42[7]^b42[6], b42[6]^b42[1], b42[0]^b42[7], b42[6]^b42[7], b42[6]};
		b43_4 = {b43[5], b43[4], b43[3]^ b43[7], b43[2]^ b43[7]^b43[6], b43[6]^b43[1], b43[0]^b43[7], b43[6]^b43[7], b43[6]};
		b44_4 = {b44[5], b44[4], b44[3]^ b44[7], b44[2]^ b44[7]^b44[6], b44[6]^b44[1], b44[0]^b44[7], b44[6]^b44[7], b44[6]};
		b45_4 = {b45[5], b45[4], b45[3]^ b45[7], b45[2]^ b45[7]^b45[6], b45[6]^b45[1], b45[0]^b45[7], b45[6]^b45[7], b45[6]};
		b46_4 = {b46[5], b46[4], b46[3]^ b46[7], b46[2]^ b46[7]^b46[6], b46[6]^b46[1], b46[0]^b46[7], b46[6]^b46[7], b46[6]};
		b47_4 = {b47[5], b47[4], b47[3]^ b47[7], b47[2]^ b47[7]^b47[6], b47[6]^b47[1], b47[0]^b47[7], b47[6]^b47[7], b47[6]};

		m4 = {
			b40_2 ^ b41_2 ^ b42_2 ^ b42 ^ b43_4 ^ b44_4 ^ b44 ^ b45_2 ^ b45 ^ b46_4 ^ b46 ^ b47_4 ^ b47_2 ^ b47,
			b41_2 ^ b42_2 ^ b43_2 ^ b43 ^ b44_4 ^ b45_4 ^ b45 ^ b46_2 ^ b46 ^ b47_4 ^ b47 ^ b40_4 ^ b40_2 ^ b40,
			b42_2 ^ b43_2 ^ b44_2 ^ b44 ^ b45_4 ^ b46_4 ^ b46 ^ b47_2 ^ b47 ^ b40_4 ^ b40 ^ b41_4 ^ b41_2 ^ b41,
			b43_2 ^ b44_2 ^ b45_2 ^ b45 ^ b46_4 ^ b47_4 ^ b47 ^ b40_2 ^ b40 ^ b41_4 ^ b41 ^ b42_4 ^ b42_2 ^ b42,
			b44_2 ^ b45_2 ^ b46_2 ^ b46 ^ b47_4 ^ b40_4 ^ b40 ^ b41_2 ^ b41 ^ b42_4 ^ b42 ^ b43_4 ^ b43_2 ^ b43,
			b45_2 ^ b46_2 ^ b47_2 ^ b47 ^ b40_4 ^ b41_4 ^ b41 ^ b42_2 ^ b42 ^ b43_4 ^ b43 ^ b44_4 ^ b44_2 ^ b44,
			b46_2 ^ b47_2 ^ b40_2 ^ b40 ^ b41_4 ^ b42_4 ^ b42 ^ b43_2 ^ b43 ^ b44_4 ^ b44 ^ b45_4 ^ b45_2 ^ b45,
			b47_2 ^ b40_2 ^ b41_2 ^ b41 ^ b42_4 ^ b43_4 ^ b43 ^ b44_2 ^ b44 ^ b45_4 ^ b45 ^ b46_4 ^ b46_2 ^ b46
		};

	end

	reg [7:0] b50,b51,b52,b53,b54,b55,b56,b57;
	reg [7:0] b50_2,b51_2,b52_2,b53_2,b54_2,b55_2,b56_2,b57_2;
	reg [7:0] b50_4,b51_4,b52_4,b53_4,b54_4,b55_4,b56_4,b57_4;

	always @ (*) begin
	
		{ b50, b51, b52, b53, b54, b55, b56, b57 } = in[703:640];
		
		b50_2 = {b50[6], b50[5], b50[4], b50[3]^b50[7], b50[2]^b50[7], b50[1], b50[0]^b50[7], b50[7]};
		b51_2 = {b51[6], b51[5], b51[4], b51[3]^b51[7], b51[2]^b51[7], b51[1], b51[0]^b51[7], b51[7]};
		b52_2 = {b52[6], b52[5], b52[4], b52[3]^b52[7], b52[2]^b52[7], b52[1], b52[0]^b52[7], b52[7]};
		b53_2 = {b53[6], b53[5], b53[4], b53[3]^b53[7], b53[2]^b53[7], b53[1], b53[0]^b53[7], b53[7]};
		b54_2 = {b54[6], b54[5], b54[4], b54[3]^b54[7], b54[2]^b54[7], b54[1], b54[0]^b54[7], b54[7]};
		b55_2 = {b55[6], b55[5], b55[4], b55[3]^b55[7], b55[2]^b55[7], b55[1], b55[0]^b55[7], b55[7]};
		b56_2 = {b56[6], b56[5], b56[4], b56[3]^b56[7], b56[2]^b56[7], b56[1], b56[0]^b56[7], b56[7]};
		b57_2 = {b57[6], b57[5], b57[4], b57[3]^b57[7], b57[2]^b57[7], b57[1], b57[0]^b57[7], b57[7]};

		b50_4 = {b50[5], b50[4], b50[3]^ b50[7], b50[2]^ b50[7]^b50[6], b50[6]^b50[1], b50[0]^b50[7], b50[6]^b50[7], b50[6]};
		b51_4 = {b51[5], b51[4], b51[3]^ b51[7], b51[2]^ b51[7]^b51[6], b51[6]^b51[1], b51[0]^b51[7], b51[6]^b51[7], b51[6]};
		b52_4 = {b52[5], b52[4], b52[3]^ b52[7], b52[2]^ b52[7]^b52[6], b52[6]^b52[1], b52[0]^b52[7], b52[6]^b52[7], b52[6]};
		b53_4 = {b53[5], b53[4], b53[3]^ b53[7], b53[2]^ b53[7]^b53[6], b53[6]^b53[1], b53[0]^b53[7], b53[6]^b53[7], b53[6]};
		b54_4 = {b54[5], b54[4], b54[3]^ b54[7], b54[2]^ b54[7]^b54[6], b54[6]^b54[1], b54[0]^b54[7], b54[6]^b54[7], b54[6]};
		b55_4 = {b55[5], b55[4], b55[3]^ b55[7], b55[2]^ b55[7]^b55[6], b55[6]^b55[1], b55[0]^b55[7], b55[6]^b55[7], b55[6]};
		b56_4 = {b56[5], b56[4], b56[3]^ b56[7], b56[2]^ b56[7]^b56[6], b56[6]^b56[1], b56[0]^b56[7], b56[6]^b56[7], b56[6]};
		b57_4 = {b57[5], b57[4], b57[3]^ b57[7], b57[2]^ b57[7]^b57[6], b57[6]^b57[1], b57[0]^b57[7], b57[6]^b57[7], b57[6]};

		m5 = {
			b50_2 ^ b51_2 ^ b52_2 ^ b52 ^ b53_4 ^ b54_4 ^ b54 ^ b55_2 ^ b55 ^ b56_4 ^ b56 ^ b57_4 ^ b57_2 ^ b57,
			b51_2 ^ b52_2 ^ b53_2 ^ b53 ^ b54_4 ^ b55_4 ^ b55 ^ b56_2 ^ b56 ^ b57_4 ^ b57 ^ b50_4 ^ b50_2 ^ b50,
			b52_2 ^ b53_2 ^ b54_2 ^ b54 ^ b55_4 ^ b56_4 ^ b56 ^ b57_2 ^ b57 ^ b50_4 ^ b50 ^ b51_4 ^ b51_2 ^ b51,
			b53_2 ^ b54_2 ^ b55_2 ^ b55 ^ b56_4 ^ b57_4 ^ b57 ^ b50_2 ^ b50 ^ b51_4 ^ b51 ^ b52_4 ^ b52_2 ^ b52,
			b54_2 ^ b55_2 ^ b56_2 ^ b56 ^ b57_4 ^ b50_4 ^ b50 ^ b51_2 ^ b51 ^ b52_4 ^ b52 ^ b53_4 ^ b53_2 ^ b53,
			b55_2 ^ b56_2 ^ b57_2 ^ b57 ^ b50_4 ^ b51_4 ^ b51 ^ b52_2 ^ b52 ^ b53_4 ^ b53 ^ b54_4 ^ b54_2 ^ b54,
			b56_2 ^ b57_2 ^ b50_2 ^ b50 ^ b51_4 ^ b52_4 ^ b52 ^ b53_2 ^ b53 ^ b54_4 ^ b54 ^ b55_4 ^ b55_2 ^ b55,
			b57_2 ^ b50_2 ^ b51_2 ^ b51 ^ b52_4 ^ b53_4 ^ b53 ^ b54_2 ^ b54 ^ b55_4 ^ b55 ^ b56_4 ^ b56_2 ^ b56
		};

	end

	reg [7:0] b60,b61,b62,b63,b64,b65,b66,b67;
	reg [7:0] b60_2,b61_2,b62_2,b63_2,b64_2,b65_2,b66_2,b67_2;
	reg [7:0] b60_4,b61_4,b62_4,b63_4,b64_4,b65_4,b66_4,b67_4;

	always @ (*) begin
	
		{ b60, b61, b62, b63, b64, b65, b66, b67 } = in[639:576];
		
		b60_2 = {b60[6], b60[5], b60[4], b60[3]^b60[7], b60[2]^b60[7], b60[1], b60[0]^b60[7], b60[7]};
		b61_2 = {b61[6], b61[5], b61[4], b61[3]^b61[7], b61[2]^b61[7], b61[1], b61[0]^b61[7], b61[7]};
		b62_2 = {b62[6], b62[5], b62[4], b62[3]^b62[7], b62[2]^b62[7], b62[1], b62[0]^b62[7], b62[7]};
		b63_2 = {b63[6], b63[5], b63[4], b63[3]^b63[7], b63[2]^b63[7], b63[1], b63[0]^b63[7], b63[7]};
		b64_2 = {b64[6], b64[5], b64[4], b64[3]^b64[7], b64[2]^b64[7], b64[1], b64[0]^b64[7], b64[7]};
		b65_2 = {b65[6], b65[5], b65[4], b65[3]^b65[7], b65[2]^b65[7], b65[1], b65[0]^b65[7], b65[7]};
		b66_2 = {b66[6], b66[5], b66[4], b66[3]^b66[7], b66[2]^b66[7], b66[1], b66[0]^b66[7], b66[7]};
		b67_2 = {b67[6], b67[5], b67[4], b67[3]^b67[7], b67[2]^b67[7], b67[1], b67[0]^b67[7], b67[7]};

		b60_4 = {b60[5], b60[4], b60[3]^ b60[7], b60[2]^ b60[7]^b60[6], b60[6]^b60[1], b60[0]^b60[7], b60[6]^b60[7], b60[6]};
		b61_4 = {b61[5], b61[4], b61[3]^ b61[7], b61[2]^ b61[7]^b61[6], b61[6]^b61[1], b61[0]^b61[7], b61[6]^b61[7], b61[6]};
		b62_4 = {b62[5], b62[4], b62[3]^ b62[7], b62[2]^ b62[7]^b62[6], b62[6]^b62[1], b62[0]^b62[7], b62[6]^b62[7], b62[6]};
		b63_4 = {b63[5], b63[4], b63[3]^ b63[7], b63[2]^ b63[7]^b63[6], b63[6]^b63[1], b63[0]^b63[7], b63[6]^b63[7], b63[6]};
		b64_4 = {b64[5], b64[4], b64[3]^ b64[7], b64[2]^ b64[7]^b64[6], b64[6]^b64[1], b64[0]^b64[7], b64[6]^b64[7], b64[6]};
		b65_4 = {b65[5], b65[4], b65[3]^ b65[7], b65[2]^ b65[7]^b65[6], b65[6]^b65[1], b65[0]^b65[7], b65[6]^b65[7], b65[6]};
		b66_4 = {b66[5], b66[4], b66[3]^ b66[7], b66[2]^ b66[7]^b66[6], b66[6]^b66[1], b66[0]^b66[7], b66[6]^b66[7], b66[6]};
		b67_4 = {b67[5], b67[4], b67[3]^ b67[7], b67[2]^ b67[7]^b67[6], b67[6]^b67[1], b67[0]^b67[7], b67[6]^b67[7], b67[6]};

		m6 = {
			b60_2 ^ b61_2 ^ b62_2 ^ b62 ^ b63_4 ^ b64_4 ^ b64 ^ b65_2 ^ b65 ^ b66_4 ^ b66 ^ b67_4 ^ b67_2 ^ b67,
			b61_2 ^ b62_2 ^ b63_2 ^ b63 ^ b64_4 ^ b65_4 ^ b65 ^ b66_2 ^ b66 ^ b67_4 ^ b67 ^ b60_4 ^ b60_2 ^ b60,
			b62_2 ^ b63_2 ^ b64_2 ^ b64 ^ b65_4 ^ b66_4 ^ b66 ^ b67_2 ^ b67 ^ b60_4 ^ b60 ^ b61_4 ^ b61_2 ^ b61,
			b63_2 ^ b64_2 ^ b65_2 ^ b65 ^ b66_4 ^ b67_4 ^ b67 ^ b60_2 ^ b60 ^ b61_4 ^ b61 ^ b62_4 ^ b62_2 ^ b62,
			b64_2 ^ b65_2 ^ b66_2 ^ b66 ^ b67_4 ^ b60_4 ^ b60 ^ b61_2 ^ b61 ^ b62_4 ^ b62 ^ b63_4 ^ b63_2 ^ b63,
			b65_2 ^ b66_2 ^ b67_2 ^ b67 ^ b60_4 ^ b61_4 ^ b61 ^ b62_2 ^ b62 ^ b63_4 ^ b63 ^ b64_4 ^ b64_2 ^ b64,
			b66_2 ^ b67_2 ^ b60_2 ^ b60 ^ b61_4 ^ b62_4 ^ b62 ^ b63_2 ^ b63 ^ b64_4 ^ b64 ^ b65_4 ^ b65_2 ^ b65,
			b67_2 ^ b60_2 ^ b61_2 ^ b61 ^ b62_4 ^ b63_4 ^ b63 ^ b64_2 ^ b64 ^ b65_4 ^ b65 ^ b66_4 ^ b66_2 ^ b66
		};

	end

	reg [7:0] b70,b71,b72,b73,b74,b75,b76,b77;
	reg [7:0] b70_2,b71_2,b72_2,b73_2,b74_2,b75_2,b76_2,b77_2;
	reg [7:0] b70_4,b71_4,b72_4,b73_4,b74_4,b75_4,b76_4,b77_4;

	always @ (*) begin
	
		{ b70, b71, b72, b73, b74, b75, b76, b77 } = in[575:512];
		
		b70_2 = {b70[6], b70[5], b70[4], b70[3]^b70[7], b70[2]^b70[7], b70[1], b70[0]^b70[7], b70[7]};
		b71_2 = {b71[6], b71[5], b71[4], b71[3]^b71[7], b71[2]^b71[7], b71[1], b71[0]^b71[7], b71[7]};
		b72_2 = {b72[6], b72[5], b72[4], b72[3]^b72[7], b72[2]^b72[7], b72[1], b72[0]^b72[7], b72[7]};
		b73_2 = {b73[6], b73[5], b73[4], b73[3]^b73[7], b73[2]^b73[7], b73[1], b73[0]^b73[7], b73[7]};
		b74_2 = {b74[6], b74[5], b74[4], b74[3]^b74[7], b74[2]^b74[7], b74[1], b74[0]^b74[7], b74[7]};
		b75_2 = {b75[6], b75[5], b75[4], b75[3]^b75[7], b75[2]^b75[7], b75[1], b75[0]^b75[7], b75[7]};
		b76_2 = {b76[6], b76[5], b76[4], b76[3]^b76[7], b76[2]^b76[7], b76[1], b76[0]^b76[7], b76[7]};
		b77_2 = {b77[6], b77[5], b77[4], b77[3]^b77[7], b77[2]^b77[7], b77[1], b77[0]^b77[7], b77[7]};

		b70_4 = {b70[5], b70[4], b70[3]^ b70[7], b70[2]^ b70[7]^b70[6], b70[6]^b70[1], b70[0]^b70[7], b70[6]^b70[7], b70[6]};
		b71_4 = {b71[5], b71[4], b71[3]^ b71[7], b71[2]^ b71[7]^b71[6], b71[6]^b71[1], b71[0]^b71[7], b71[6]^b71[7], b71[6]};
		b72_4 = {b72[5], b72[4], b72[3]^ b72[7], b72[2]^ b72[7]^b72[6], b72[6]^b72[1], b72[0]^b72[7], b72[6]^b72[7], b72[6]};
		b73_4 = {b73[5], b73[4], b73[3]^ b73[7], b73[2]^ b73[7]^b73[6], b73[6]^b73[1], b73[0]^b73[7], b73[6]^b73[7], b73[6]};
		b74_4 = {b74[5], b74[4], b74[3]^ b74[7], b74[2]^ b74[7]^b74[6], b74[6]^b74[1], b74[0]^b74[7], b74[6]^b74[7], b74[6]};
		b75_4 = {b75[5], b75[4], b75[3]^ b75[7], b75[2]^ b75[7]^b75[6], b75[6]^b75[1], b75[0]^b75[7], b75[6]^b75[7], b75[6]};
		b76_4 = {b76[5], b76[4], b76[3]^ b76[7], b76[2]^ b76[7]^b76[6], b76[6]^b76[1], b76[0]^b76[7], b76[6]^b76[7], b76[6]};
		b77_4 = {b77[5], b77[4], b77[3]^ b77[7], b77[2]^ b77[7]^b77[6], b77[6]^b77[1], b77[0]^b77[7], b77[6]^b77[7], b77[6]};

		m7 = {
			b70_2 ^ b71_2 ^ b72_2 ^ b72 ^ b73_4 ^ b74_4 ^ b74 ^ b75_2 ^ b75 ^ b76_4 ^ b76 ^ b77_4 ^ b77_2 ^ b77,
			b71_2 ^ b72_2 ^ b73_2 ^ b73 ^ b74_4 ^ b75_4 ^ b75 ^ b76_2 ^ b76 ^ b77_4 ^ b77 ^ b70_4 ^ b70_2 ^ b70,
			b72_2 ^ b73_2 ^ b74_2 ^ b74 ^ b75_4 ^ b76_4 ^ b76 ^ b77_2 ^ b77 ^ b70_4 ^ b70 ^ b71_4 ^ b71_2 ^ b71,
			b73_2 ^ b74_2 ^ b75_2 ^ b75 ^ b76_4 ^ b77_4 ^ b77 ^ b70_2 ^ b70 ^ b71_4 ^ b71 ^ b72_4 ^ b72_2 ^ b72,
			b74_2 ^ b75_2 ^ b76_2 ^ b76 ^ b77_4 ^ b70_4 ^ b70 ^ b71_2 ^ b71 ^ b72_4 ^ b72 ^ b73_4 ^ b73_2 ^ b73,
			b75_2 ^ b76_2 ^ b77_2 ^ b77 ^ b70_4 ^ b71_4 ^ b71 ^ b72_2 ^ b72 ^ b73_4 ^ b73 ^ b74_4 ^ b74_2 ^ b74,
			b76_2 ^ b77_2 ^ b70_2 ^ b70 ^ b71_4 ^ b72_4 ^ b72 ^ b73_2 ^ b73 ^ b74_4 ^ b74 ^ b75_4 ^ b75_2 ^ b75,
			b77_2 ^ b70_2 ^ b71_2 ^ b71 ^ b72_4 ^ b73_4 ^ b73 ^ b74_2 ^ b74 ^ b75_4 ^ b75 ^ b76_4 ^ b76_2 ^ b76
		};

	end

	reg [7:0] b80,b81,b82,b83,b84,b85,b86,b87;
	reg [7:0] b80_2,b81_2,b82_2,b83_2,b84_2,b85_2,b86_2,b87_2;
	reg [7:0] b80_4,b81_4,b82_4,b83_4,b84_4,b85_4,b86_4,b87_4;

	always @ (*) begin
	
		{ b80, b81, b82, b83, b84, b85, b86, b87 } = in[511:448];
		
		b80_2 = {b80[6], b80[5], b80[4], b80[3]^b80[7], b80[2]^b80[7], b80[1], b80[0]^b80[7], b80[7]};
		b81_2 = {b81[6], b81[5], b81[4], b81[3]^b81[7], b81[2]^b81[7], b81[1], b81[0]^b81[7], b81[7]};
		b82_2 = {b82[6], b82[5], b82[4], b82[3]^b82[7], b82[2]^b82[7], b82[1], b82[0]^b82[7], b82[7]};
		b83_2 = {b83[6], b83[5], b83[4], b83[3]^b83[7], b83[2]^b83[7], b83[1], b83[0]^b83[7], b83[7]};
		b84_2 = {b84[6], b84[5], b84[4], b84[3]^b84[7], b84[2]^b84[7], b84[1], b84[0]^b84[7], b84[7]};
		b85_2 = {b85[6], b85[5], b85[4], b85[3]^b85[7], b85[2]^b85[7], b85[1], b85[0]^b85[7], b85[7]};
		b86_2 = {b86[6], b86[5], b86[4], b86[3]^b86[7], b86[2]^b86[7], b86[1], b86[0]^b86[7], b86[7]};
		b87_2 = {b87[6], b87[5], b87[4], b87[3]^b87[7], b87[2]^b87[7], b87[1], b87[0]^b87[7], b87[7]};

		b80_4 = {b80[5], b80[4], b80[3]^ b80[7], b80[2]^ b80[7]^b80[6], b80[6]^b80[1], b80[0]^b80[7], b80[6]^b80[7], b80[6]};
		b81_4 = {b81[5], b81[4], b81[3]^ b81[7], b81[2]^ b81[7]^b81[6], b81[6]^b81[1], b81[0]^b81[7], b81[6]^b81[7], b81[6]};
		b82_4 = {b82[5], b82[4], b82[3]^ b82[7], b82[2]^ b82[7]^b82[6], b82[6]^b82[1], b82[0]^b82[7], b82[6]^b82[7], b82[6]};
		b83_4 = {b83[5], b83[4], b83[3]^ b83[7], b83[2]^ b83[7]^b83[6], b83[6]^b83[1], b83[0]^b83[7], b83[6]^b83[7], b83[6]};
		b84_4 = {b84[5], b84[4], b84[3]^ b84[7], b84[2]^ b84[7]^b84[6], b84[6]^b84[1], b84[0]^b84[7], b84[6]^b84[7], b84[6]};
		b85_4 = {b85[5], b85[4], b85[3]^ b85[7], b85[2]^ b85[7]^b85[6], b85[6]^b85[1], b85[0]^b85[7], b85[6]^b85[7], b85[6]};
		b86_4 = {b86[5], b86[4], b86[3]^ b86[7], b86[2]^ b86[7]^b86[6], b86[6]^b86[1], b86[0]^b86[7], b86[6]^b86[7], b86[6]};
		b87_4 = {b87[5], b87[4], b87[3]^ b87[7], b87[2]^ b87[7]^b87[6], b87[6]^b87[1], b87[0]^b87[7], b87[6]^b87[7], b87[6]};

		m8 = {
			b80_2 ^ b81_2 ^ b82_2 ^ b82 ^ b83_4 ^ b84_4 ^ b84 ^ b85_2 ^ b85 ^ b86_4 ^ b86 ^ b87_4 ^ b87_2 ^ b87,
			b81_2 ^ b82_2 ^ b83_2 ^ b83 ^ b84_4 ^ b85_4 ^ b85 ^ b86_2 ^ b86 ^ b87_4 ^ b87 ^ b80_4 ^ b80_2 ^ b80,
			b82_2 ^ b83_2 ^ b84_2 ^ b84 ^ b85_4 ^ b86_4 ^ b86 ^ b87_2 ^ b87 ^ b80_4 ^ b80 ^ b81_4 ^ b81_2 ^ b81,
			b83_2 ^ b84_2 ^ b85_2 ^ b85 ^ b86_4 ^ b87_4 ^ b87 ^ b80_2 ^ b80 ^ b81_4 ^ b81 ^ b82_4 ^ b82_2 ^ b82,
			b84_2 ^ b85_2 ^ b86_2 ^ b86 ^ b87_4 ^ b80_4 ^ b80 ^ b81_2 ^ b81 ^ b82_4 ^ b82 ^ b83_4 ^ b83_2 ^ b83,
			b85_2 ^ b86_2 ^ b87_2 ^ b87 ^ b80_4 ^ b81_4 ^ b81 ^ b82_2 ^ b82 ^ b83_4 ^ b83 ^ b84_4 ^ b84_2 ^ b84,
			b86_2 ^ b87_2 ^ b80_2 ^ b80 ^ b81_4 ^ b82_4 ^ b82 ^ b83_2 ^ b83 ^ b84_4 ^ b84 ^ b85_4 ^ b85_2 ^ b85,
			b87_2 ^ b80_2 ^ b81_2 ^ b81 ^ b82_4 ^ b83_4 ^ b83 ^ b84_2 ^ b84 ^ b85_4 ^ b85 ^ b86_4 ^ b86_2 ^ b86
		};

	end

	reg [7:0] b90,b91,b92,b93,b94,b95,b96,b97;
	reg [7:0] b90_2,b91_2,b92_2,b93_2,b94_2,b95_2,b96_2,b97_2;
	reg [7:0] b90_4,b91_4,b92_4,b93_4,b94_4,b95_4,b96_4,b97_4;

	always @ (*) begin
	
		{ b90, b91, b92, b93, b94, b95, b96, b97 } = in[447:384];
		
		b90_2 = {b90[6], b90[5], b90[4], b90[3]^b90[7], b90[2]^b90[7], b90[1], b90[0]^b90[7], b90[7]};
		b91_2 = {b91[6], b91[5], b91[4], b91[3]^b91[7], b91[2]^b91[7], b91[1], b91[0]^b91[7], b91[7]};
		b92_2 = {b92[6], b92[5], b92[4], b92[3]^b92[7], b92[2]^b92[7], b92[1], b92[0]^b92[7], b92[7]};
		b93_2 = {b93[6], b93[5], b93[4], b93[3]^b93[7], b93[2]^b93[7], b93[1], b93[0]^b93[7], b93[7]};
		b94_2 = {b94[6], b94[5], b94[4], b94[3]^b94[7], b94[2]^b94[7], b94[1], b94[0]^b94[7], b94[7]};
		b95_2 = {b95[6], b95[5], b95[4], b95[3]^b95[7], b95[2]^b95[7], b95[1], b95[0]^b95[7], b95[7]};
		b96_2 = {b96[6], b96[5], b96[4], b96[3]^b96[7], b96[2]^b96[7], b96[1], b96[0]^b96[7], b96[7]};
		b97_2 = {b97[6], b97[5], b97[4], b97[3]^b97[7], b97[2]^b97[7], b97[1], b97[0]^b97[7], b97[7]};

		b90_4 = {b90[5], b90[4], b90[3]^ b90[7], b90[2]^ b90[7]^b90[6], b90[6]^b90[1], b90[0]^b90[7], b90[6]^b90[7], b90[6]};
		b91_4 = {b91[5], b91[4], b91[3]^ b91[7], b91[2]^ b91[7]^b91[6], b91[6]^b91[1], b91[0]^b91[7], b91[6]^b91[7], b91[6]};
		b92_4 = {b92[5], b92[4], b92[3]^ b92[7], b92[2]^ b92[7]^b92[6], b92[6]^b92[1], b92[0]^b92[7], b92[6]^b92[7], b92[6]};
		b93_4 = {b93[5], b93[4], b93[3]^ b93[7], b93[2]^ b93[7]^b93[6], b93[6]^b93[1], b93[0]^b93[7], b93[6]^b93[7], b93[6]};
		b94_4 = {b94[5], b94[4], b94[3]^ b94[7], b94[2]^ b94[7]^b94[6], b94[6]^b94[1], b94[0]^b94[7], b94[6]^b94[7], b94[6]};
		b95_4 = {b95[5], b95[4], b95[3]^ b95[7], b95[2]^ b95[7]^b95[6], b95[6]^b95[1], b95[0]^b95[7], b95[6]^b95[7], b95[6]};
		b96_4 = {b96[5], b96[4], b96[3]^ b96[7], b96[2]^ b96[7]^b96[6], b96[6]^b96[1], b96[0]^b96[7], b96[6]^b96[7], b96[6]};
		b97_4 = {b97[5], b97[4], b97[3]^ b97[7], b97[2]^ b97[7]^b97[6], b97[6]^b97[1], b97[0]^b97[7], b97[6]^b97[7], b97[6]};

		m9 = {
			b90_2 ^ b91_2 ^ b92_2 ^ b92 ^ b93_4 ^ b94_4 ^ b94 ^ b95_2 ^ b95 ^ b96_4 ^ b96 ^ b97_4 ^ b97_2 ^ b97,
			b91_2 ^ b92_2 ^ b93_2 ^ b93 ^ b94_4 ^ b95_4 ^ b95 ^ b96_2 ^ b96 ^ b97_4 ^ b97 ^ b90_4 ^ b90_2 ^ b90,
			b92_2 ^ b93_2 ^ b94_2 ^ b94 ^ b95_4 ^ b96_4 ^ b96 ^ b97_2 ^ b97 ^ b90_4 ^ b90 ^ b91_4 ^ b91_2 ^ b91,
			b93_2 ^ b94_2 ^ b95_2 ^ b95 ^ b96_4 ^ b97_4 ^ b97 ^ b90_2 ^ b90 ^ b91_4 ^ b91 ^ b92_4 ^ b92_2 ^ b92,
			b94_2 ^ b95_2 ^ b96_2 ^ b96 ^ b97_4 ^ b90_4 ^ b90 ^ b91_2 ^ b91 ^ b92_4 ^ b92 ^ b93_4 ^ b93_2 ^ b93,
			b95_2 ^ b96_2 ^ b97_2 ^ b97 ^ b90_4 ^ b91_4 ^ b91 ^ b92_2 ^ b92 ^ b93_4 ^ b93 ^ b94_4 ^ b94_2 ^ b94,
			b96_2 ^ b97_2 ^ b90_2 ^ b90 ^ b91_4 ^ b92_4 ^ b92 ^ b93_2 ^ b93 ^ b94_4 ^ b94 ^ b95_4 ^ b95_2 ^ b95,
			b97_2 ^ b90_2 ^ b91_2 ^ b91 ^ b92_4 ^ b93_4 ^ b93 ^ b94_2 ^ b94 ^ b95_4 ^ b95 ^ b96_4 ^ b96_2 ^ b96
		};

	end

	reg [7:0] bA0,bA1,bA2,bA3,bA4,bA5,bA6,bA7;
	reg [7:0] bA0_2,bA1_2,bA2_2,bA3_2,bA4_2,bA5_2,bA6_2,bA7_2;
	reg [7:0] bA0_4,bA1_4,bA2_4,bA3_4,bA4_4,bA5_4,bA6_4,bA7_4;

	always @ (*) begin
	
		{ bA0, bA1, bA2, bA3, bA4, bA5, bA6, bA7 } = in[383:320];
		
		bA0_2 = {bA0[6], bA0[5], bA0[4], bA0[3]^bA0[7], bA0[2]^bA0[7], bA0[1], bA0[0]^bA0[7], bA0[7]};
		bA1_2 = {bA1[6], bA1[5], bA1[4], bA1[3]^bA1[7], bA1[2]^bA1[7], bA1[1], bA1[0]^bA1[7], bA1[7]};
		bA2_2 = {bA2[6], bA2[5], bA2[4], bA2[3]^bA2[7], bA2[2]^bA2[7], bA2[1], bA2[0]^bA2[7], bA2[7]};
		bA3_2 = {bA3[6], bA3[5], bA3[4], bA3[3]^bA3[7], bA3[2]^bA3[7], bA3[1], bA3[0]^bA3[7], bA3[7]};
		bA4_2 = {bA4[6], bA4[5], bA4[4], bA4[3]^bA4[7], bA4[2]^bA4[7], bA4[1], bA4[0]^bA4[7], bA4[7]};
		bA5_2 = {bA5[6], bA5[5], bA5[4], bA5[3]^bA5[7], bA5[2]^bA5[7], bA5[1], bA5[0]^bA5[7], bA5[7]};
		bA6_2 = {bA6[6], bA6[5], bA6[4], bA6[3]^bA6[7], bA6[2]^bA6[7], bA6[1], bA6[0]^bA6[7], bA6[7]};
		bA7_2 = {bA7[6], bA7[5], bA7[4], bA7[3]^bA7[7], bA7[2]^bA7[7], bA7[1], bA7[0]^bA7[7], bA7[7]};

		bA0_4 = {bA0[5], bA0[4], bA0[3]^ bA0[7], bA0[2]^ bA0[7]^bA0[6], bA0[6]^bA0[1], bA0[0]^bA0[7], bA0[6]^bA0[7], bA0[6]};
		bA1_4 = {bA1[5], bA1[4], bA1[3]^ bA1[7], bA1[2]^ bA1[7]^bA1[6], bA1[6]^bA1[1], bA1[0]^bA1[7], bA1[6]^bA1[7], bA1[6]};
		bA2_4 = {bA2[5], bA2[4], bA2[3]^ bA2[7], bA2[2]^ bA2[7]^bA2[6], bA2[6]^bA2[1], bA2[0]^bA2[7], bA2[6]^bA2[7], bA2[6]};
		bA3_4 = {bA3[5], bA3[4], bA3[3]^ bA3[7], bA3[2]^ bA3[7]^bA3[6], bA3[6]^bA3[1], bA3[0]^bA3[7], bA3[6]^bA3[7], bA3[6]};
		bA4_4 = {bA4[5], bA4[4], bA4[3]^ bA4[7], bA4[2]^ bA4[7]^bA4[6], bA4[6]^bA4[1], bA4[0]^bA4[7], bA4[6]^bA4[7], bA4[6]};
		bA5_4 = {bA5[5], bA5[4], bA5[3]^ bA5[7], bA5[2]^ bA5[7]^bA5[6], bA5[6]^bA5[1], bA5[0]^bA5[7], bA5[6]^bA5[7], bA5[6]};
		bA6_4 = {bA6[5], bA6[4], bA6[3]^ bA6[7], bA6[2]^ bA6[7]^bA6[6], bA6[6]^bA6[1], bA6[0]^bA6[7], bA6[6]^bA6[7], bA6[6]};
		bA7_4 = {bA7[5], bA7[4], bA7[3]^ bA7[7], bA7[2]^ bA7[7]^bA7[6], bA7[6]^bA7[1], bA7[0]^bA7[7], bA7[6]^bA7[7], bA7[6]};

		mA = {
			bA0_2 ^ bA1_2 ^ bA2_2 ^ bA2 ^ bA3_4 ^ bA4_4 ^ bA4 ^ bA5_2 ^ bA5 ^ bA6_4 ^ bA6 ^ bA7_4 ^ bA7_2 ^ bA7,
			bA1_2 ^ bA2_2 ^ bA3_2 ^ bA3 ^ bA4_4 ^ bA5_4 ^ bA5 ^ bA6_2 ^ bA6 ^ bA7_4 ^ bA7 ^ bA0_4 ^ bA0_2 ^ bA0,
			bA2_2 ^ bA3_2 ^ bA4_2 ^ bA4 ^ bA5_4 ^ bA6_4 ^ bA6 ^ bA7_2 ^ bA7 ^ bA0_4 ^ bA0 ^ bA1_4 ^ bA1_2 ^ bA1,
			bA3_2 ^ bA4_2 ^ bA5_2 ^ bA5 ^ bA6_4 ^ bA7_4 ^ bA7 ^ bA0_2 ^ bA0 ^ bA1_4 ^ bA1 ^ bA2_4 ^ bA2_2 ^ bA2,
			bA4_2 ^ bA5_2 ^ bA6_2 ^ bA6 ^ bA7_4 ^ bA0_4 ^ bA0 ^ bA1_2 ^ bA1 ^ bA2_4 ^ bA2 ^ bA3_4 ^ bA3_2 ^ bA3,
			bA5_2 ^ bA6_2 ^ bA7_2 ^ bA7 ^ bA0_4 ^ bA1_4 ^ bA1 ^ bA2_2 ^ bA2 ^ bA3_4 ^ bA3 ^ bA4_4 ^ bA4_2 ^ bA4,
			bA6_2 ^ bA7_2 ^ bA0_2 ^ bA0 ^ bA1_4 ^ bA2_4 ^ bA2 ^ bA3_2 ^ bA3 ^ bA4_4 ^ bA4 ^ bA5_4 ^ bA5_2 ^ bA5,
			bA7_2 ^ bA0_2 ^ bA1_2 ^ bA1 ^ bA2_4 ^ bA3_4 ^ bA3 ^ bA4_2 ^ bA4 ^ bA5_4 ^ bA5 ^ bA6_4 ^ bA6_2 ^ bA6
		};

	end

	reg [7:0] bB0,bB1,bB2,bB3,bB4,bB5,bB6,bB7;
	reg [7:0] bB0_2,bB1_2,bB2_2,bB3_2,bB4_2,bB5_2,bB6_2,bB7_2;
	reg [7:0] bB0_4,bB1_4,bB2_4,bB3_4,bB4_4,bB5_4,bB6_4,bB7_4;

	always @ (*) begin
	
		{ bB0, bB1, bB2, bB3, bB4, bB5, bB6, bB7 } = in[319:256];
		
		bB0_2 = {bB0[6], bB0[5], bB0[4], bB0[3]^bB0[7], bB0[2]^bB0[7], bB0[1], bB0[0]^bB0[7], bB0[7]};
		bB1_2 = {bB1[6], bB1[5], bB1[4], bB1[3]^bB1[7], bB1[2]^bB1[7], bB1[1], bB1[0]^bB1[7], bB1[7]};
		bB2_2 = {bB2[6], bB2[5], bB2[4], bB2[3]^bB2[7], bB2[2]^bB2[7], bB2[1], bB2[0]^bB2[7], bB2[7]};
		bB3_2 = {bB3[6], bB3[5], bB3[4], bB3[3]^bB3[7], bB3[2]^bB3[7], bB3[1], bB3[0]^bB3[7], bB3[7]};
		bB4_2 = {bB4[6], bB4[5], bB4[4], bB4[3]^bB4[7], bB4[2]^bB4[7], bB4[1], bB4[0]^bB4[7], bB4[7]};
		bB5_2 = {bB5[6], bB5[5], bB5[4], bB5[3]^bB5[7], bB5[2]^bB5[7], bB5[1], bB5[0]^bB5[7], bB5[7]};
		bB6_2 = {bB6[6], bB6[5], bB6[4], bB6[3]^bB6[7], bB6[2]^bB6[7], bB6[1], bB6[0]^bB6[7], bB6[7]};
		bB7_2 = {bB7[6], bB7[5], bB7[4], bB7[3]^bB7[7], bB7[2]^bB7[7], bB7[1], bB7[0]^bB7[7], bB7[7]};

		bB0_4 = {bB0[5], bB0[4], bB0[3]^ bB0[7], bB0[2]^ bB0[7]^bB0[6], bB0[6]^bB0[1], bB0[0]^bB0[7], bB0[6]^bB0[7], bB0[6]};
		bB1_4 = {bB1[5], bB1[4], bB1[3]^ bB1[7], bB1[2]^ bB1[7]^bB1[6], bB1[6]^bB1[1], bB1[0]^bB1[7], bB1[6]^bB1[7], bB1[6]};
		bB2_4 = {bB2[5], bB2[4], bB2[3]^ bB2[7], bB2[2]^ bB2[7]^bB2[6], bB2[6]^bB2[1], bB2[0]^bB2[7], bB2[6]^bB2[7], bB2[6]};
		bB3_4 = {bB3[5], bB3[4], bB3[3]^ bB3[7], bB3[2]^ bB3[7]^bB3[6], bB3[6]^bB3[1], bB3[0]^bB3[7], bB3[6]^bB3[7], bB3[6]};
		bB4_4 = {bB4[5], bB4[4], bB4[3]^ bB4[7], bB4[2]^ bB4[7]^bB4[6], bB4[6]^bB4[1], bB4[0]^bB4[7], bB4[6]^bB4[7], bB4[6]};
		bB5_4 = {bB5[5], bB5[4], bB5[3]^ bB5[7], bB5[2]^ bB5[7]^bB5[6], bB5[6]^bB5[1], bB5[0]^bB5[7], bB5[6]^bB5[7], bB5[6]};
		bB6_4 = {bB6[5], bB6[4], bB6[3]^ bB6[7], bB6[2]^ bB6[7]^bB6[6], bB6[6]^bB6[1], bB6[0]^bB6[7], bB6[6]^bB6[7], bB6[6]};
		bB7_4 = {bB7[5], bB7[4], bB7[3]^ bB7[7], bB7[2]^ bB7[7]^bB7[6], bB7[6]^bB7[1], bB7[0]^bB7[7], bB7[6]^bB7[7], bB7[6]};

		mB = {
			bB0_2 ^ bB1_2 ^ bB2_2 ^ bB2 ^ bB3_4 ^ bB4_4 ^ bB4 ^ bB5_2 ^ bB5 ^ bB6_4 ^ bB6 ^ bB7_4 ^ bB7_2 ^ bB7,
			bB1_2 ^ bB2_2 ^ bB3_2 ^ bB3 ^ bB4_4 ^ bB5_4 ^ bB5 ^ bB6_2 ^ bB6 ^ bB7_4 ^ bB7 ^ bB0_4 ^ bB0_2 ^ bB0,
			bB2_2 ^ bB3_2 ^ bB4_2 ^ bB4 ^ bB5_4 ^ bB6_4 ^ bB6 ^ bB7_2 ^ bB7 ^ bB0_4 ^ bB0 ^ bB1_4 ^ bB1_2 ^ bB1,
			bB3_2 ^ bB4_2 ^ bB5_2 ^ bB5 ^ bB6_4 ^ bB7_4 ^ bB7 ^ bB0_2 ^ bB0 ^ bB1_4 ^ bB1 ^ bB2_4 ^ bB2_2 ^ bB2,
			bB4_2 ^ bB5_2 ^ bB6_2 ^ bB6 ^ bB7_4 ^ bB0_4 ^ bB0 ^ bB1_2 ^ bB1 ^ bB2_4 ^ bB2 ^ bB3_4 ^ bB3_2 ^ bB3,
			bB5_2 ^ bB6_2 ^ bB7_2 ^ bB7 ^ bB0_4 ^ bB1_4 ^ bB1 ^ bB2_2 ^ bB2 ^ bB3_4 ^ bB3 ^ bB4_4 ^ bB4_2 ^ bB4,
			bB6_2 ^ bB7_2 ^ bB0_2 ^ bB0 ^ bB1_4 ^ bB2_4 ^ bB2 ^ bB3_2 ^ bB3 ^ bB4_4 ^ bB4 ^ bB5_4 ^ bB5_2 ^ bB5,
			bB7_2 ^ bB0_2 ^ bB1_2 ^ bB1 ^ bB2_4 ^ bB3_4 ^ bB3 ^ bB4_2 ^ bB4 ^ bB5_4 ^ bB5 ^ bB6_4 ^ bB6_2 ^ bB6
		};

	end

	reg [7:0] bC0,bC1,bC2,bC3,bC4,bC5,bC6,bC7;
	reg [7:0] bC0_2,bC1_2,bC2_2,bC3_2,bC4_2,bC5_2,bC6_2,bC7_2;
	reg [7:0] bC0_4,bC1_4,bC2_4,bC3_4,bC4_4,bC5_4,bC6_4,bC7_4;

	always @ (*) begin
	
		{ bC0, bC1, bC2, bC3, bC4, bC5, bC6, bC7 } = in[255:192];
		
		bC0_2 = {bC0[6], bC0[5], bC0[4], bC0[3]^bC0[7], bC0[2]^bC0[7], bC0[1], bC0[0]^bC0[7], bC0[7]};
		bC1_2 = {bC1[6], bC1[5], bC1[4], bC1[3]^bC1[7], bC1[2]^bC1[7], bC1[1], bC1[0]^bC1[7], bC1[7]};
		bC2_2 = {bC2[6], bC2[5], bC2[4], bC2[3]^bC2[7], bC2[2]^bC2[7], bC2[1], bC2[0]^bC2[7], bC2[7]};
		bC3_2 = {bC3[6], bC3[5], bC3[4], bC3[3]^bC3[7], bC3[2]^bC3[7], bC3[1], bC3[0]^bC3[7], bC3[7]};
		bC4_2 = {bC4[6], bC4[5], bC4[4], bC4[3]^bC4[7], bC4[2]^bC4[7], bC4[1], bC4[0]^bC4[7], bC4[7]};
		bC5_2 = {bC5[6], bC5[5], bC5[4], bC5[3]^bC5[7], bC5[2]^bC5[7], bC5[1], bC5[0]^bC5[7], bC5[7]};
		bC6_2 = {bC6[6], bC6[5], bC6[4], bC6[3]^bC6[7], bC6[2]^bC6[7], bC6[1], bC6[0]^bC6[7], bC6[7]};
		bC7_2 = {bC7[6], bC7[5], bC7[4], bC7[3]^bC7[7], bC7[2]^bC7[7], bC7[1], bC7[0]^bC7[7], bC7[7]};

		bC0_4 = {bC0[5], bC0[4], bC0[3]^ bC0[7], bC0[2]^ bC0[7]^bC0[6], bC0[6]^bC0[1], bC0[0]^bC0[7], bC0[6]^bC0[7], bC0[6]};
		bC1_4 = {bC1[5], bC1[4], bC1[3]^ bC1[7], bC1[2]^ bC1[7]^bC1[6], bC1[6]^bC1[1], bC1[0]^bC1[7], bC1[6]^bC1[7], bC1[6]};
		bC2_4 = {bC2[5], bC2[4], bC2[3]^ bC2[7], bC2[2]^ bC2[7]^bC2[6], bC2[6]^bC2[1], bC2[0]^bC2[7], bC2[6]^bC2[7], bC2[6]};
		bC3_4 = {bC3[5], bC3[4], bC3[3]^ bC3[7], bC3[2]^ bC3[7]^bC3[6], bC3[6]^bC3[1], bC3[0]^bC3[7], bC3[6]^bC3[7], bC3[6]};
		bC4_4 = {bC4[5], bC4[4], bC4[3]^ bC4[7], bC4[2]^ bC4[7]^bC4[6], bC4[6]^bC4[1], bC4[0]^bC4[7], bC4[6]^bC4[7], bC4[6]};
		bC5_4 = {bC5[5], bC5[4], bC5[3]^ bC5[7], bC5[2]^ bC5[7]^bC5[6], bC5[6]^bC5[1], bC5[0]^bC5[7], bC5[6]^bC5[7], bC5[6]};
		bC6_4 = {bC6[5], bC6[4], bC6[3]^ bC6[7], bC6[2]^ bC6[7]^bC6[6], bC6[6]^bC6[1], bC6[0]^bC6[7], bC6[6]^bC6[7], bC6[6]};
		bC7_4 = {bC7[5], bC7[4], bC7[3]^ bC7[7], bC7[2]^ bC7[7]^bC7[6], bC7[6]^bC7[1], bC7[0]^bC7[7], bC7[6]^bC7[7], bC7[6]};

		mC = {
			bC0_2 ^ bC1_2 ^ bC2_2 ^ bC2 ^ bC3_4 ^ bC4_4 ^ bC4 ^ bC5_2 ^ bC5 ^ bC6_4 ^ bC6 ^ bC7_4 ^ bC7_2 ^ bC7,
			bC1_2 ^ bC2_2 ^ bC3_2 ^ bC3 ^ bC4_4 ^ bC5_4 ^ bC5 ^ bC6_2 ^ bC6 ^ bC7_4 ^ bC7 ^ bC0_4 ^ bC0_2 ^ bC0,
			bC2_2 ^ bC3_2 ^ bC4_2 ^ bC4 ^ bC5_4 ^ bC6_4 ^ bC6 ^ bC7_2 ^ bC7 ^ bC0_4 ^ bC0 ^ bC1_4 ^ bC1_2 ^ bC1,
			bC3_2 ^ bC4_2 ^ bC5_2 ^ bC5 ^ bC6_4 ^ bC7_4 ^ bC7 ^ bC0_2 ^ bC0 ^ bC1_4 ^ bC1 ^ bC2_4 ^ bC2_2 ^ bC2,
			bC4_2 ^ bC5_2 ^ bC6_2 ^ bC6 ^ bC7_4 ^ bC0_4 ^ bC0 ^ bC1_2 ^ bC1 ^ bC2_4 ^ bC2 ^ bC3_4 ^ bC3_2 ^ bC3,
			bC5_2 ^ bC6_2 ^ bC7_2 ^ bC7 ^ bC0_4 ^ bC1_4 ^ bC1 ^ bC2_2 ^ bC2 ^ bC3_4 ^ bC3 ^ bC4_4 ^ bC4_2 ^ bC4,
			bC6_2 ^ bC7_2 ^ bC0_2 ^ bC0 ^ bC1_4 ^ bC2_4 ^ bC2 ^ bC3_2 ^ bC3 ^ bC4_4 ^ bC4 ^ bC5_4 ^ bC5_2 ^ bC5,
			bC7_2 ^ bC0_2 ^ bC1_2 ^ bC1 ^ bC2_4 ^ bC3_4 ^ bC3 ^ bC4_2 ^ bC4 ^ bC5_4 ^ bC5 ^ bC6_4 ^ bC6_2 ^ bC6
		};

	end

	reg [7:0] bD0,bD1,bD2,bD3,bD4,bD5,bD6,bD7;
	reg [7:0] bD0_2,bD1_2,bD2_2,bD3_2,bD4_2,bD5_2,bD6_2,bD7_2;
	reg [7:0] bD0_4,bD1_4,bD2_4,bD3_4,bD4_4,bD5_4,bD6_4,bD7_4;

	always @ (*) begin
	
		{ bD0, bD1, bD2, bD3, bD4, bD5, bD6, bD7 } = in[191:128];
		
		bD0_2 = {bD0[6], bD0[5], bD0[4], bD0[3]^bD0[7], bD0[2]^bD0[7], bD0[1], bD0[0]^bD0[7], bD0[7]};
		bD1_2 = {bD1[6], bD1[5], bD1[4], bD1[3]^bD1[7], bD1[2]^bD1[7], bD1[1], bD1[0]^bD1[7], bD1[7]};
		bD2_2 = {bD2[6], bD2[5], bD2[4], bD2[3]^bD2[7], bD2[2]^bD2[7], bD2[1], bD2[0]^bD2[7], bD2[7]};
		bD3_2 = {bD3[6], bD3[5], bD3[4], bD3[3]^bD3[7], bD3[2]^bD3[7], bD3[1], bD3[0]^bD3[7], bD3[7]};
		bD4_2 = {bD4[6], bD4[5], bD4[4], bD4[3]^bD4[7], bD4[2]^bD4[7], bD4[1], bD4[0]^bD4[7], bD4[7]};
		bD5_2 = {bD5[6], bD5[5], bD5[4], bD5[3]^bD5[7], bD5[2]^bD5[7], bD5[1], bD5[0]^bD5[7], bD5[7]};
		bD6_2 = {bD6[6], bD6[5], bD6[4], bD6[3]^bD6[7], bD6[2]^bD6[7], bD6[1], bD6[0]^bD6[7], bD6[7]};
		bD7_2 = {bD7[6], bD7[5], bD7[4], bD7[3]^bD7[7], bD7[2]^bD7[7], bD7[1], bD7[0]^bD7[7], bD7[7]};

		bD0_4 = {bD0[5], bD0[4], bD0[3]^ bD0[7], bD0[2]^ bD0[7]^bD0[6], bD0[6]^bD0[1], bD0[0]^bD0[7], bD0[6]^bD0[7], bD0[6]};
		bD1_4 = {bD1[5], bD1[4], bD1[3]^ bD1[7], bD1[2]^ bD1[7]^bD1[6], bD1[6]^bD1[1], bD1[0]^bD1[7], bD1[6]^bD1[7], bD1[6]};
		bD2_4 = {bD2[5], bD2[4], bD2[3]^ bD2[7], bD2[2]^ bD2[7]^bD2[6], bD2[6]^bD2[1], bD2[0]^bD2[7], bD2[6]^bD2[7], bD2[6]};
		bD3_4 = {bD3[5], bD3[4], bD3[3]^ bD3[7], bD3[2]^ bD3[7]^bD3[6], bD3[6]^bD3[1], bD3[0]^bD3[7], bD3[6]^bD3[7], bD3[6]};
		bD4_4 = {bD4[5], bD4[4], bD4[3]^ bD4[7], bD4[2]^ bD4[7]^bD4[6], bD4[6]^bD4[1], bD4[0]^bD4[7], bD4[6]^bD4[7], bD4[6]};
		bD5_4 = {bD5[5], bD5[4], bD5[3]^ bD5[7], bD5[2]^ bD5[7]^bD5[6], bD5[6]^bD5[1], bD5[0]^bD5[7], bD5[6]^bD5[7], bD5[6]};
		bD6_4 = {bD6[5], bD6[4], bD6[3]^ bD6[7], bD6[2]^ bD6[7]^bD6[6], bD6[6]^bD6[1], bD6[0]^bD6[7], bD6[6]^bD6[7], bD6[6]};
		bD7_4 = {bD7[5], bD7[4], bD7[3]^ bD7[7], bD7[2]^ bD7[7]^bD7[6], bD7[6]^bD7[1], bD7[0]^bD7[7], bD7[6]^bD7[7], bD7[6]};

		mD = {
			bD0_2 ^ bD1_2 ^ bD2_2 ^ bD2 ^ bD3_4 ^ bD4_4 ^ bD4 ^ bD5_2 ^ bD5 ^ bD6_4 ^ bD6 ^ bD7_4 ^ bD7_2 ^ bD7,
			bD1_2 ^ bD2_2 ^ bD3_2 ^ bD3 ^ bD4_4 ^ bD5_4 ^ bD5 ^ bD6_2 ^ bD6 ^ bD7_4 ^ bD7 ^ bD0_4 ^ bD0_2 ^ bD0,
			bD2_2 ^ bD3_2 ^ bD4_2 ^ bD4 ^ bD5_4 ^ bD6_4 ^ bD6 ^ bD7_2 ^ bD7 ^ bD0_4 ^ bD0 ^ bD1_4 ^ bD1_2 ^ bD1,
			bD3_2 ^ bD4_2 ^ bD5_2 ^ bD5 ^ bD6_4 ^ bD7_4 ^ bD7 ^ bD0_2 ^ bD0 ^ bD1_4 ^ bD1 ^ bD2_4 ^ bD2_2 ^ bD2,
			bD4_2 ^ bD5_2 ^ bD6_2 ^ bD6 ^ bD7_4 ^ bD0_4 ^ bD0 ^ bD1_2 ^ bD1 ^ bD2_4 ^ bD2 ^ bD3_4 ^ bD3_2 ^ bD3,
			bD5_2 ^ bD6_2 ^ bD7_2 ^ bD7 ^ bD0_4 ^ bD1_4 ^ bD1 ^ bD2_2 ^ bD2 ^ bD3_4 ^ bD3 ^ bD4_4 ^ bD4_2 ^ bD4,
			bD6_2 ^ bD7_2 ^ bD0_2 ^ bD0 ^ bD1_4 ^ bD2_4 ^ bD2 ^ bD3_2 ^ bD3 ^ bD4_4 ^ bD4 ^ bD5_4 ^ bD5_2 ^ bD5,
			bD7_2 ^ bD0_2 ^ bD1_2 ^ bD1 ^ bD2_4 ^ bD3_4 ^ bD3 ^ bD4_2 ^ bD4 ^ bD5_4 ^ bD5 ^ bD6_4 ^ bD6_2 ^ bD6
		};

	end

	reg [7:0] bE0,bE1,bE2,bE3,bE4,bE5,bE6,bE7;
	reg [7:0] bE0_2,bE1_2,bE2_2,bE3_2,bE4_2,bE5_2,bE6_2,bE7_2;
	reg [7:0] bE0_4,bE1_4,bE2_4,bE3_4,bE4_4,bE5_4,bE6_4,bE7_4;

	always @ (*) begin
	
		{ bE0, bE1, bE2, bE3, bE4, bE5, bE6, bE7 } = in[127:64];
		
		bE0_2 = {bE0[6], bE0[5], bE0[4], bE0[3]^bE0[7], bE0[2]^bE0[7], bE0[1], bE0[0]^bE0[7], bE0[7]};
		bE1_2 = {bE1[6], bE1[5], bE1[4], bE1[3]^bE1[7], bE1[2]^bE1[7], bE1[1], bE1[0]^bE1[7], bE1[7]};
		bE2_2 = {bE2[6], bE2[5], bE2[4], bE2[3]^bE2[7], bE2[2]^bE2[7], bE2[1], bE2[0]^bE2[7], bE2[7]};
		bE3_2 = {bE3[6], bE3[5], bE3[4], bE3[3]^bE3[7], bE3[2]^bE3[7], bE3[1], bE3[0]^bE3[7], bE3[7]};
		bE4_2 = {bE4[6], bE4[5], bE4[4], bE4[3]^bE4[7], bE4[2]^bE4[7], bE4[1], bE4[0]^bE4[7], bE4[7]};
		bE5_2 = {bE5[6], bE5[5], bE5[4], bE5[3]^bE5[7], bE5[2]^bE5[7], bE5[1], bE5[0]^bE5[7], bE5[7]};
		bE6_2 = {bE6[6], bE6[5], bE6[4], bE6[3]^bE6[7], bE6[2]^bE6[7], bE6[1], bE6[0]^bE6[7], bE6[7]};
		bE7_2 = {bE7[6], bE7[5], bE7[4], bE7[3]^bE7[7], bE7[2]^bE7[7], bE7[1], bE7[0]^bE7[7], bE7[7]};

		bE0_4 = {bE0[5], bE0[4], bE0[3]^ bE0[7], bE0[2]^ bE0[7]^bE0[6], bE0[6]^bE0[1], bE0[0]^bE0[7], bE0[6]^bE0[7], bE0[6]};
		bE1_4 = {bE1[5], bE1[4], bE1[3]^ bE1[7], bE1[2]^ bE1[7]^bE1[6], bE1[6]^bE1[1], bE1[0]^bE1[7], bE1[6]^bE1[7], bE1[6]};
		bE2_4 = {bE2[5], bE2[4], bE2[3]^ bE2[7], bE2[2]^ bE2[7]^bE2[6], bE2[6]^bE2[1], bE2[0]^bE2[7], bE2[6]^bE2[7], bE2[6]};
		bE3_4 = {bE3[5], bE3[4], bE3[3]^ bE3[7], bE3[2]^ bE3[7]^bE3[6], bE3[6]^bE3[1], bE3[0]^bE3[7], bE3[6]^bE3[7], bE3[6]};
		bE4_4 = {bE4[5], bE4[4], bE4[3]^ bE4[7], bE4[2]^ bE4[7]^bE4[6], bE4[6]^bE4[1], bE4[0]^bE4[7], bE4[6]^bE4[7], bE4[6]};
		bE5_4 = {bE5[5], bE5[4], bE5[3]^ bE5[7], bE5[2]^ bE5[7]^bE5[6], bE5[6]^bE5[1], bE5[0]^bE5[7], bE5[6]^bE5[7], bE5[6]};
		bE6_4 = {bE6[5], bE6[4], bE6[3]^ bE6[7], bE6[2]^ bE6[7]^bE6[6], bE6[6]^bE6[1], bE6[0]^bE6[7], bE6[6]^bE6[7], bE6[6]};
		bE7_4 = {bE7[5], bE7[4], bE7[3]^ bE7[7], bE7[2]^ bE7[7]^bE7[6], bE7[6]^bE7[1], bE7[0]^bE7[7], bE7[6]^bE7[7], bE7[6]};

		mE = {
			bE0_2 ^ bE1_2 ^ bE2_2 ^ bE2 ^ bE3_4 ^ bE4_4 ^ bE4 ^ bE5_2 ^ bE5 ^ bE6_4 ^ bE6 ^ bE7_4 ^ bE7_2 ^ bE7,
			bE1_2 ^ bE2_2 ^ bE3_2 ^ bE3 ^ bE4_4 ^ bE5_4 ^ bE5 ^ bE6_2 ^ bE6 ^ bE7_4 ^ bE7 ^ bE0_4 ^ bE0_2 ^ bE0,
			bE2_2 ^ bE3_2 ^ bE4_2 ^ bE4 ^ bE5_4 ^ bE6_4 ^ bE6 ^ bE7_2 ^ bE7 ^ bE0_4 ^ bE0 ^ bE1_4 ^ bE1_2 ^ bE1,
			bE3_2 ^ bE4_2 ^ bE5_2 ^ bE5 ^ bE6_4 ^ bE7_4 ^ bE7 ^ bE0_2 ^ bE0 ^ bE1_4 ^ bE1 ^ bE2_4 ^ bE2_2 ^ bE2,
			bE4_2 ^ bE5_2 ^ bE6_2 ^ bE6 ^ bE7_4 ^ bE0_4 ^ bE0 ^ bE1_2 ^ bE1 ^ bE2_4 ^ bE2 ^ bE3_4 ^ bE3_2 ^ bE3,
			bE5_2 ^ bE6_2 ^ bE7_2 ^ bE7 ^ bE0_4 ^ bE1_4 ^ bE1 ^ bE2_2 ^ bE2 ^ bE3_4 ^ bE3 ^ bE4_4 ^ bE4_2 ^ bE4,
			bE6_2 ^ bE7_2 ^ bE0_2 ^ bE0 ^ bE1_4 ^ bE2_4 ^ bE2 ^ bE3_2 ^ bE3 ^ bE4_4 ^ bE4 ^ bE5_4 ^ bE5_2 ^ bE5,
			bE7_2 ^ bE0_2 ^ bE1_2 ^ bE1 ^ bE2_4 ^ bE3_4 ^ bE3 ^ bE4_2 ^ bE4 ^ bE5_4 ^ bE5 ^ bE6_4 ^ bE6_2 ^ bE6
		};

	end

	reg [7:0] bF0,bF1,bF2,bF3,bF4,bF5,bF6,bF7;
	reg [7:0] bF0_2,bF1_2,bF2_2,bF3_2,bF4_2,bF5_2,bF6_2,bF7_2;
	reg [7:0] bF0_4,bF1_4,bF2_4,bF3_4,bF4_4,bF5_4,bF6_4,bF7_4;

	always @ (*) begin
	
		{ bF0, bF1, bF2, bF3, bF4, bF5, bF6, bF7 } = in[63:0];
		
		bF0_2 = {bF0[6], bF0[5], bF0[4], bF0[3]^bF0[7], bF0[2]^bF0[7], bF0[1], bF0[0]^bF0[7], bF0[7]};
		bF1_2 = {bF1[6], bF1[5], bF1[4], bF1[3]^bF1[7], bF1[2]^bF1[7], bF1[1], bF1[0]^bF1[7], bF1[7]};
		bF2_2 = {bF2[6], bF2[5], bF2[4], bF2[3]^bF2[7], bF2[2]^bF2[7], bF2[1], bF2[0]^bF2[7], bF2[7]};
		bF3_2 = {bF3[6], bF3[5], bF3[4], bF3[3]^bF3[7], bF3[2]^bF3[7], bF3[1], bF3[0]^bF3[7], bF3[7]};
		bF4_2 = {bF4[6], bF4[5], bF4[4], bF4[3]^bF4[7], bF4[2]^bF4[7], bF4[1], bF4[0]^bF4[7], bF4[7]};
		bF5_2 = {bF5[6], bF5[5], bF5[4], bF5[3]^bF5[7], bF5[2]^bF5[7], bF5[1], bF5[0]^bF5[7], bF5[7]};
		bF6_2 = {bF6[6], bF6[5], bF6[4], bF6[3]^bF6[7], bF6[2]^bF6[7], bF6[1], bF6[0]^bF6[7], bF6[7]};
		bF7_2 = {bF7[6], bF7[5], bF7[4], bF7[3]^bF7[7], bF7[2]^bF7[7], bF7[1], bF7[0]^bF7[7], bF7[7]};

		bF0_4 = {bF0[5], bF0[4], bF0[3]^ bF0[7], bF0[2]^ bF0[7]^bF0[6], bF0[6]^bF0[1], bF0[0]^bF0[7], bF0[6]^bF0[7], bF0[6]};
		bF1_4 = {bF1[5], bF1[4], bF1[3]^ bF1[7], bF1[2]^ bF1[7]^bF1[6], bF1[6]^bF1[1], bF1[0]^bF1[7], bF1[6]^bF1[7], bF1[6]};
		bF2_4 = {bF2[5], bF2[4], bF2[3]^ bF2[7], bF2[2]^ bF2[7]^bF2[6], bF2[6]^bF2[1], bF2[0]^bF2[7], bF2[6]^bF2[7], bF2[6]};
		bF3_4 = {bF3[5], bF3[4], bF3[3]^ bF3[7], bF3[2]^ bF3[7]^bF3[6], bF3[6]^bF3[1], bF3[0]^bF3[7], bF3[6]^bF3[7], bF3[6]};
		bF4_4 = {bF4[5], bF4[4], bF4[3]^ bF4[7], bF4[2]^ bF4[7]^bF4[6], bF4[6]^bF4[1], bF4[0]^bF4[7], bF4[6]^bF4[7], bF4[6]};
		bF5_4 = {bF5[5], bF5[4], bF5[3]^ bF5[7], bF5[2]^ bF5[7]^bF5[6], bF5[6]^bF5[1], bF5[0]^bF5[7], bF5[6]^bF5[7], bF5[6]};
		bF6_4 = {bF6[5], bF6[4], bF6[3]^ bF6[7], bF6[2]^ bF6[7]^bF6[6], bF6[6]^bF6[1], bF6[0]^bF6[7], bF6[6]^bF6[7], bF6[6]};
		bF7_4 = {bF7[5], bF7[4], bF7[3]^ bF7[7], bF7[2]^ bF7[7]^bF7[6], bF7[6]^bF7[1], bF7[0]^bF7[7], bF7[6]^bF7[7], bF7[6]};

		mF = {
			bF0_2 ^ bF1_2 ^ bF2_2 ^ bF2 ^ bF3_4 ^ bF4_4 ^ bF4 ^ bF5_2 ^ bF5 ^ bF6_4 ^ bF6 ^ bF7_4 ^ bF7_2 ^ bF7,
			bF1_2 ^ bF2_2 ^ bF3_2 ^ bF3 ^ bF4_4 ^ bF5_4 ^ bF5 ^ bF6_2 ^ bF6 ^ bF7_4 ^ bF7 ^ bF0_4 ^ bF0_2 ^ bF0,
			bF2_2 ^ bF3_2 ^ bF4_2 ^ bF4 ^ bF5_4 ^ bF6_4 ^ bF6 ^ bF7_2 ^ bF7 ^ bF0_4 ^ bF0 ^ bF1_4 ^ bF1_2 ^ bF1,
			bF3_2 ^ bF4_2 ^ bF5_2 ^ bF5 ^ bF6_4 ^ bF7_4 ^ bF7 ^ bF0_2 ^ bF0 ^ bF1_4 ^ bF1 ^ bF2_4 ^ bF2_2 ^ bF2,
			bF4_2 ^ bF5_2 ^ bF6_2 ^ bF6 ^ bF7_4 ^ bF0_4 ^ bF0 ^ bF1_2 ^ bF1 ^ bF2_4 ^ bF2 ^ bF3_4 ^ bF3_2 ^ bF3,
			bF5_2 ^ bF6_2 ^ bF7_2 ^ bF7 ^ bF0_4 ^ bF1_4 ^ bF1 ^ bF2_2 ^ bF2 ^ bF3_4 ^ bF3 ^ bF4_4 ^ bF4_2 ^ bF4,
			bF6_2 ^ bF7_2 ^ bF0_2 ^ bF0 ^ bF1_4 ^ bF2_4 ^ bF2 ^ bF3_2 ^ bF3 ^ bF4_4 ^ bF4 ^ bF5_4 ^ bF5_2 ^ bF5,
			bF7_2 ^ bF0_2 ^ bF1_2 ^ bF1 ^ bF2_4 ^ bF3_4 ^ bF3 ^ bF4_2 ^ bF4 ^ bF5_4 ^ bF5 ^ bF6_4 ^ bF6_2 ^ bF6
		};

	end

	always @ (posedge clk) begin
		out <= {m0,m1,m2,m3,m4,m5,m6,m7,m8,m9,mA,mB,mC,mD,mE,mF};
	end

endmodule
