/*
 * Copyright (c) 2017 Sprocket
 *
 * This is free software: you can redistribute it and/or modify
 * it under the terms of the GNU Affero General Public License with
 * additional permissions to the one published by the Free Software
 * Foundation, either version 3 of the License, or (at your option)
 * any later version. For more information see LICENSE.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU Affero General Public License for more details.
 *
 * You should have received a copy of the GNU Affero General Public License
 * along with this program. If not, see <http://www.gnu.org/licenses/>.
 */

module fugue512 (
	input clk,
	input [511:0] data,
	output [511:0] hash
);

	reg [511:0] H;
	assign hash = H;

	reg [511:0] x0, x0_1, x0_2, x0_3, x0_4, x0_5, x0_6, x0_7;
	reg [479:0] x1, x1_1, x1_2, x1_3, x1_4, x1_5, x1_6, x1_7, x1_8;
	reg [447:0] x2, x2_1, x2_2, x2_3, x2_4, x2_5, x2_6, x2_7, x2_8;
	reg [415:0] x3, x3_1, x3_2, x3_3, x3_4, x3_5, x3_6, x3_7, x3_8;
	reg [383:0] x4, x4_1, x4_2, x4_3, x4_4, x4_5, x4_6, x4_7, x4_8;
	reg [351:0] x5, x5_1, x5_2, x5_3, x5_4, x5_5, x5_6, x5_7, x5_8;
	reg [319:0] x6, x6_1, x6_2, x6_3, x6_4, x6_5, x6_6, x6_7, x6_8;
	reg [287:0] x7, x7_1, x7_2, x7_3, x7_4, x7_5, x7_6, x7_7, x7_8;
	reg [255:0] x8, x8_1, x8_2, x8_3, x8_4, x8_5, x8_6, x8_7, x8_8;
	reg [223:0] x9, x9_1, x9_2, x9_3, x9_4, x9_5, x9_6, x9_7, x9_8;
	reg [191:0] x10, x10_1, x10_2, x10_3, x10_4, x10_5, x10_6, x10_7, x10_8;
	reg [159:0] x11, x11_1, x11_2, x11_3, x11_4, x11_5, x11_6, x11_7, x11_8;
	reg [127:0] x12, x12_1, x12_2, x12_3, x12_4, x12_5, x12_6, x12_7, x12_8;
	reg [ 95:0] x13, x13_1, x13_2, x13_3, x13_4, x13_5, x13_6, x13_7, x13_8;
	reg [ 63:0] x14, x14_1, x14_2, x14_3, x14_4, x14_5, x14_6, x14_7, x14_8;
	reg [ 31:0] x15, x15_1, x15_2, x15_3, x15_4, x15_5, x15_6, x15_7, x15_8;
	
	reg [1151:0] S0;

	wire [1151:0] S1,S2,S3,S4,S5,S6,S7,S8,S9,S10,S11,S12,S13,S14,S15,S16,S17,S18;
	wire [1151:0] C0,C1,C2,C3,C4,C5,C6,C7,C8,C9,C10,C11,C12,C13,C14,C15;
	wire [1151:0] C16,C17,C18,C19,C20,C21,C22,C23,C24,C25,C26,C27,C28,C29,C30,C31,C32;	
	wire [1151:0] D0,D1,D2,D3,D4,D5,D6,D7,D8,D9,D10,D11,D12;
	
	round r0  (clk, x0[511:480], S0,  S1);
	round r1  (clk, x1[479:448], S1,  S2);
	round r2  (clk, x2[447:416], S2,  S3);
	round r3  (clk, x3[415:384], S3,  S4);
	round r4  (clk, x4[383:352], S4,  S5);
	round r5  (clk, x5[351:320], S5,  S6);
	round r6  (clk, x6[319:288], S6,  S7);
	round r7  (clk, x7[287:256], S7,  S8);
	round r8  (clk, x8[255:224], S8,  S9);
	round r9  (clk, x9[223:192], S9,  S10);
	round r10 (clk, x10[191:160], S10, S11);
	round r11 (clk, x11[159:128], S11, S12);
	round r12 (clk, x12[127: 96], S12, S13);
	round r13 (clk, x13[ 95: 64], S13, S14);
	round r14 (clk, x14[ 63: 32], S14, S15);
	round r15 (clk, x15[ 31:  0], S15, S16);
	round r16 (clk, 32'h00000000,  S16, S17);
	round r17 (clk, 32'h00000200,  S17, S18);
	
	close_1 c0 (clk, { S18[1055:0], S18[1151:1056] }, C0);
	close_1 c1 (clk, C0, C1);
	close_1 c2 (clk, C1, C2);
	close_1 c3 (clk, C2, C3);
	close_1 c4 (clk, C3, C4);
	close_1 c5 (clk, C4, C5);
	close_1 c6 (clk, C5, C6);
	close_1 c7 (clk, C6, C7);
	close_1 c8 (clk, C7, C8);
	close_1 c9 (clk, C8, C9);
	close_1 c10 (clk, C9, C10);
	close_1 c11 (clk, C10, C11);
	close_1 c12 (clk, C11, C12);
	close_1 c13 (clk, C12, C13);
	close_1 c14 (clk, C13, C14);
	close_1 c15 (clk, C14, C15);
	close_1 c16 (clk, C15, C16);
	close_1 c17 (clk, C16, C17);
	close_1 c18 (clk, C17, C18);
	close_1 c19 (clk, C18, C19);
	close_1 c20 (clk, C19, C20);
	close_1 c21 (clk, C20, C21);
	close_1 c22 (clk, C21, C22);
	close_1 c23 (clk, C22, C23);
	close_1 c24 (clk, C23, C24);
	close_1 c25 (clk, C24, C25);
	close_1 c26 (clk, C25, C26);
	close_1 c27 (clk, C26, C27);
	close_1 c28 (clk, C27, C28);
	close_1 c29 (clk, C28, C29);
	close_1 c30 (clk, C29, C30);
	close_1 c31 (clk, C30, C31);

	close_2 d0 (clk, { C31[95:0], C31[1151:96] }, D0);
	close_2 d1 (clk, D0, D1);
	close_2 d2 (clk, D1, D2);
	close_2 d3 (clk, D2, D3);
	close_2 d4 (clk, D3, D4);
	close_2 d5 (clk, D4, D5);
	close_2 d6 (clk, D5, D6);
	close_2 d7 (clk, D6, D7);
	close_2 d8 (clk, D7, D8);
	close_2 d9 (clk, D8, D9);
	close_2 d10 (clk, D9, D10);
	close_2 d11 (clk, D10, D11);
	close_2 d12 (clk, D11, D12);
	
	always @ (posedge clk) begin

		S0[1151:640] <= 512'he13e3567da6ed11d951fddd625ea78e7437f203fcae65838ddb21398aac6e2c94a92efd106e8020bb6eecc54d915f117ac9ab027c5d3e4dbe616af758807a57e;
		S0[639:0] <= 640'd0;
	
		x15 = x15_7;
		x15_8 = x15_7;
		x15_7 = x15_6;
		x15_6 = x15_5;
		x15_5 = x15_4;
		x15_4 = x15_3;
		x15_3 = x15_2;
		x15_2 = x15_1;
		x15_1 = x14[31:0];
		x14 = x14_7;
		x14_8 = x14_7;
		x14_7 = x14_6;
		x14_6 = x14_5;
		x14_5 = x14_4;
		x14_4 = x14_3;
		x14_3 = x14_2;
		x14_2 = x14_1;
		x14_1 = x13[63:0];
		x13 = x13_7;
		x13_8 = x13_7;
		x13_7 = x13_6;
		x13_6 = x13_5;
		x13_5 = x13_4;
		x13_4 = x13_3;
		x13_3 = x13_2;
		x13_2 = x13_1;
		x13_1 = x12[95:0];
		x12 = x12_7;
		x12_8 = x12_7;
		x12_7 = x12_6;
		x12_6 = x12_5;
		x12_5 = x12_4;
		x12_4 = x12_3;
		x12_3 = x12_2;
		x12_2 = x12_1;
		x12_1 = x11[127:0];
		x11 = x11_7;
		x11_8 = x11_7;
		x11_7 = x11_6;
		x11_6 = x11_5;
		x11_5 = x11_4;
		x11_4 = x11_3;
		x11_3 = x11_2;
		x11_2 = x11_1;
		x11_1 = x10[159:0];
		x10 = x10_7;
		x10_8 = x10_7;
		x10_7 = x10_6;
		x10_6 = x10_5;
		x10_5 = x10_4;
		x10_4 = x10_3;
		x10_3 = x10_2;
		x10_2 = x10_1;
		x10_1 = x9[191:0];
		x9 = x9_7;
		x9_8 = x9_7;
		x9_7 = x9_6;
		x9_6 = x9_5;
		x9_5 = x9_4;
		x9_4 = x9_3;
		x9_3 = x9_2;
		x9_2 = x9_1;
		x9_1 = x8[223:0];
		x8 = x8_7;
		x8_8 = x8_7;
		x8_7 = x8_6;
		x8_6 = x8_5;
		x8_5 = x8_4;
		x8_4 = x8_3;
		x8_3 = x8_2;
		x8_2 = x8_1;
		x8_1 = x7[255:0];
		x7 = x7_7;
		x7_8 = x7_7;
		x7_7 = x7_6;
		x7_6 = x7_5;
		x7_5 = x7_4;
		x7_4 = x7_3;
		x7_3 = x7_2;
		x7_2 = x7_1;
		x7_1 = x6[287:0];
		x6 = x6_7;
		x6_8 = x6_7;
		x6_7 = x6_6;
		x6_6 = x6_5;
		x6_5 = x6_4;
		x6_4 = x6_3;
		x6_3 = x6_2;
		x6_2 = x6_1;
		x6_1 = x5[319:0];
		x5 = x5_7;
		x5_8 = x5_7;
		x5_7 = x5_6;
		x5_6 = x5_5;
		x5_5 = x5_4;
		x5_4 = x5_3;
		x5_3 = x5_2;
		x5_2 = x5_1;
		x5_1 = x4[351:0];
		x4 = x4_7;
		x4_8 = x4_7;
		x4_7 = x4_6;
		x4_6 = x4_5;
		x4_5 = x4_4;
		x4_4 = x4_3;
		x4_3 = x4_2;
		x4_2 = x4_1;
		x4_1 = x3[383:0];
		x3 = x3_7;
		x3_8 = x3_7;
		x3_7 = x3_6;
		x3_6 = x3_5;
		x3_5 = x3_4;
		x3_4 = x3_3;
		x3_3 = x3_2;
		x3_2 = x3_1;
		x3_1 = x2[415:0];
		x2 = x2_7;
		x2_8 = x2_7;
		x2_7 = x2_6;
		x2_6 = x2_5;
		x2_5 = x2_4;
		x2_4 = x2_3;
		x2_3 = x2_2;
		x2_2 = x2_1;
		x2_1 = x1[447:0];
		x1 = x1_7;
		x1_8 = x1_7;
		x1_7 = x1_6;
		x1_6 = x1_5;
		x1_5 = x1_4;
		x1_4 = x1_3;
		x1_3 = x1_2;
		x1_2 = x1_1;
		x1_1 = x0[479:0];
		x0 = data;
//		x0_6 = x0_5;
//		x0_5 = x0_4;
//		x0_4 = x0_3;
//		x0_3 = x0_2;
//		x0_2 = x0_1;
//		x0_1 = data;

		H = {
			D12[ 32 +: 32],
			D12[ 64 +: 32],
			D12[ 96 +: 32],
			D12[128 +: 32] ^ D12[0 +: 32],
			D12[288 +: 32] ^ D12[0 +: 32],
			D12[320 +: 32],
			D12[352 +: 32],
			D12[384 +: 32],
			D12[576 +: 32] ^ D12[0 +: 32],
			D12[608 +: 32],
			D12[640 +: 32],
			D12[672 +: 32],
			D12[864 +: 32] ^ D12[0 +: 32],
			D12[896 +: 32],
			D12[928 +: 32],
			D12[960 +: 32]
		};
		
	end

endmodule

//module TIX (
//	input [1151:0] in,
//	input [31:0] q,
//	output [1151:0] out
//);
//
//	assign out[1152-((36- 0)*32) +: 32] = q;
//	assign out[1152-((36- 1)*32) +: 32] = in[1152-((36- 1)*32) +: 32] ^ in[1152-((36-24)*32) +: 32];
//	assign out[1152-((36- 2)*32) +: 32] = in[1152-((36- 2)*32) +: 32];
//	assign out[1152-((36- 3)*32) +: 32] = in[1152-((36- 3)*32) +: 32];
//	assign out[1152-((36- 4)*32) +: 32] = in[1152-((36- 4)*32) +: 32] ^ in[1152-((36-27)*32) +: 32];
//	assign out[1152-((36- 5)*32) +: 32] = in[1152-((36- 5)*32) +: 32];
//	assign out[1152-((36- 6)*32) +: 32] = in[1152-((36- 6)*32) +: 32];
//	assign out[1152-((36- 7)*32) +: 32] = in[1152-((36- 7)*32) +: 32] ^ in[1152-((36-30)*32) +: 32];
//	assign out[1152-((36- 8)*32) +: 32] = in[1152-((36- 8)*32) +: 32] ^ q;
//	assign out[1152-((36- 9)*32) +: 32] = in[1152-((36- 9)*32) +: 32];
//	assign out[1152-((36-10)*32) +: 32] = in[1152-((36-10)*32) +: 32];
//	assign out[1152-((36-11)*32) +: 32] = in[1152-((36-11)*32) +: 32];
//	assign out[1152-((36-12)*32) +: 32] = in[1152-((36-12)*32) +: 32];
//	assign out[1152-((36-13)*32) +: 32] = in[1152-((36-13)*32) +: 32];
//	assign out[1152-((36-14)*32) +: 32] = in[1152-((36-14)*32) +: 32];
//	assign out[1152-((36-15)*32) +: 32] = in[1152-((36-15)*32) +: 32];
//	assign out[1152-((36-16)*32) +: 32] = in[1152-((36-16)*32) +: 32];
//	assign out[1152-((36-17)*32) +: 32] = in[1152-((36-17)*32) +: 32];
//	assign out[1152-((36-18)*32) +: 32] = in[1152-((36-18)*32) +: 32];
//	assign out[1152-((36-19)*32) +: 32] = in[1152-((36-19)*32) +: 32];
//	assign out[1152-((36-20)*32) +: 32] = in[1152-((36-20)*32) +: 32];
//	assign out[1152-((36-21)*32) +: 32] = in[1152-((36-21)*32) +: 32];
//	assign out[1152-((36-22)*32) +: 32] = in[1152-((36-22)*32) +: 32] ^ in[1152-((36- 0)*32) +: 32];
//	assign out[1152-((36-23)*32) +: 32] = in[1152-((36-23)*32) +: 32];
//	assign out[1152-((36-24)*32) +: 32] = in[1152-((36-24)*32) +: 32];
//	assign out[1152-((36-25)*32) +: 32] = in[1152-((36-25)*32) +: 32];
//	assign out[1152-((36-26)*32) +: 32] = in[1152-((36-26)*32) +: 32];
//	assign out[1152-((36-27)*32) +: 32] = in[1152-((36-27)*32) +: 32];
//	assign out[1152-((36-28)*32) +: 32] = in[1152-((36-28)*32) +: 32];
//	assign out[1152-((36-29)*32) +: 32] = in[1152-((36-29)*32) +: 32];
//	assign out[1152-((36-30)*32) +: 32] = in[1152-((36-30)*32) +: 32];
//	assign out[1152-((36-31)*32) +: 32] = in[1152-((36-31)*32) +: 32];
//	assign out[1152-((36-32)*32) +: 32] = in[1152-((36-32)*32) +: 32];
//	assign out[1152-((36-33)*32) +: 32] = in[1152-((36-33)*32) +: 32];
//	assign out[1152-((36-34)*32) +: 32] = in[1152-((36-34)*32) +: 32];
//	assign out[1152-((36-35)*32) +: 32] = in[1152-((36-35)*32) +: 32];
//
//endmodule


//module CMIX (
//	input [95:0] i0,
//	input [95:0] i1,
//	input [95:0] i2,
//	output [95:0] o1,
//	output [95:0] o2
//);
//
//	assign o1 = i0 ^ i2;
//	assign o2 = i1 ^ i2;
//
//endmodule


module round (
	input clk,
	input [31:0] q,
	input [1151:0] S,
	output [1151:0] O
);

	wire [127:0] S1, S2, S3, S4;
	wire [1151:0] tix;

	wire [1151:0] S0i, S1i, S2i, S3i, S4i;
	reg [1151:0] S0ix, S1ix, S2ix, S3ix;
	reg [1151:0] S0ixx, S1ixx, S2ixx, S3ixx;

	assign tix[1152-((36- 0)*32) +: 32] = q;
	assign tix[1152-((36- 1)*32) +: 32] = S[1152-((36- 1)*32) +: 32] ^ S[1152-((36-24)*32) +: 32];
	assign tix[1152-((36- 2)*32) +: 32] = S[1152-((36- 2)*32) +: 32];
	assign tix[1152-((36- 3)*32) +: 32] = S[1152-((36- 3)*32) +: 32];
	assign tix[1152-((36- 4)*32) +: 32] = S[1152-((36- 4)*32) +: 32] ^ S[1152-((36-27)*32) +: 32];
	assign tix[1152-((36- 5)*32) +: 32] = S[1152-((36- 5)*32) +: 32];
	assign tix[1152-((36- 6)*32) +: 32] = S[1152-((36- 6)*32) +: 32];
	assign tix[1152-((36- 7)*32) +: 32] = S[1152-((36- 7)*32) +: 32] ^ S[1152-((36-30)*32) +: 32];
	assign tix[1152-((36- 8)*32) +: 32] = S[1152-((36- 8)*32) +: 32] ^ q;
	assign tix[1152-((36- 9)*32) +: 32] = S[1152-((36- 9)*32) +: 32];
	assign tix[1152-((36-10)*32) +: 32] = S[1152-((36-10)*32) +: 32];
	assign tix[1152-((36-11)*32) +: 32] = S[1152-((36-11)*32) +: 32];
	assign tix[1152-((36-12)*32) +: 32] = S[1152-((36-12)*32) +: 32];
	assign tix[1152-((36-13)*32) +: 32] = S[1152-((36-13)*32) +: 32];
	assign tix[1152-((36-14)*32) +: 32] = S[1152-((36-14)*32) +: 32];
	assign tix[1152-((36-15)*32) +: 32] = S[1152-((36-15)*32) +: 32];
	assign tix[1152-((36-16)*32) +: 32] = S[1152-((36-16)*32) +: 32];
	assign tix[1152-((36-17)*32) +: 32] = S[1152-((36-17)*32) +: 32];
	assign tix[1152-((36-18)*32) +: 32] = S[1152-((36-18)*32) +: 32];
	assign tix[1152-((36-19)*32) +: 32] = S[1152-((36-19)*32) +: 32];
	assign tix[1152-((36-20)*32) +: 32] = S[1152-((36-20)*32) +: 32];
	assign tix[1152-((36-21)*32) +: 32] = S[1152-((36-21)*32) +: 32];
	assign tix[1152-((36-22)*32) +: 32] = S[1152-((36-22)*32) +: 32] ^ S[1152-((36- 0)*32) +: 32];
	assign tix[1152-((36-23)*32) +: 32] = S[1152-((36-23)*32) +: 32];
	assign tix[1152-((36-24)*32) +: 32] = S[1152-((36-24)*32) +: 32];
	assign tix[1152-((36-25)*32) +: 32] = S[1152-((36-25)*32) +: 32];
	assign tix[1152-((36-26)*32) +: 32] = S[1152-((36-26)*32) +: 32];
	assign tix[1152-((36-27)*32) +: 32] = S[1152-((36-27)*32) +: 32];
	assign tix[1152-((36-28)*32) +: 32] = S[1152-((36-28)*32) +: 32];
	assign tix[1152-((36-29)*32) +: 32] = S[1152-((36-29)*32) +: 32];
	assign tix[1152-((36-30)*32) +: 32] = S[1152-((36-30)*32) +: 32];
	assign tix[1152-((36-31)*32) +: 32] = S[1152-((36-31)*32) +: 32];
	assign tix[1152-((36-32)*32) +: 32] = S[1152-((36-32)*32) +: 32];
	assign tix[1152-((36-33)*32) +: 32] = S[1152-((36-33)*32) +: 32];
	assign tix[1152-((36-34)*32) +: 32] = S[1152-((36-34)*32) +: 32];
	assign tix[1152-((36-35)*32) +: 32] = S[1152-((36-35)*32) +: 32];

	assign S0i[1152-((36-33)*32) +: 32] = tix[1152-((36-33)*32) +: 32] ^ tix[1152-((36- 1)*32) +: 32];
	assign S0i[1152-((36-34)*32) +: 32] = tix[1152-((36-34)*32) +: 32] ^ tix[1152-((36- 2)*32) +: 32];
	assign S0i[1152-((36-35)*32) +: 32] = tix[1152-((36-35)*32) +: 32] ^ tix[1152-((36- 3)*32) +: 32];
	assign S0i[1152-((36-15)*32) +: 32] = tix[1152-((36-15)*32) +: 32] ^ tix[1152-((36- 1)*32) +: 32];
	assign S0i[1152-((36-16)*32) +: 32] = tix[1152-((36-16)*32) +: 32] ^ tix[1152-((36- 2)*32) +: 32];
	assign S0i[1152-((36-17)*32) +: 32] = tix[1152-((36-17)*32) +: 32] ^ tix[1152-((36- 3)*32) +: 32];
	assign S0i[1151-((36-15)*32) : 1152-((36-0)*32)] = tix[1151-((36-15)*32) : 1152-((36-0)*32)];
	assign S0i[1151-((36-33)*32) : 1152-((36-18)*32)] = tix[1151-((36-33)*32) : 1152-((36-18)*32)];
	
	assign S1i[1152-((36-33)*32) +: 32] = S1[127:96];
	assign S1i[1152-((36-34)*32) +: 32] = S1[95:64];
	assign S1i[1152-((36-35)*32) +: 32] = S1[63:32];
	assign S1i[1152-((36- 0)*32) +: 32] = S1[31:0];
	assign S1i[1152-((36-30)*32) +: 32] = S0ix[1152-((36-30)*32) +: 32] ^ S1[95:64];
	assign S1i[1152-((36-31)*32) +: 32] = S0ix[1152-((36-31)*32) +: 32] ^ S1[63:32];
	assign S1i[1152-((36-32)*32) +: 32] = S0ix[1152-((36-32)*32) +: 32] ^ S1[31:0];
	assign S1i[1152-((36-12)*32) +: 32] = S0ix[1152-((36-12)*32) +: 32] ^ S1[95:64];
	assign S1i[1152-((36-13)*32) +: 32] = S0ix[1152-((36-13)*32) +: 32] ^ S1[63:32];
	assign S1i[1152-((36-14)*32) +: 32] = S0ix[1152-((36-14)*32) +: 32] ^ S1[31:0];
	assign S1i[1151-((36-12)*32) : 1152-((36-1)*32)] = S0ix[1151-((36-12)*32) : 1152-((36-1)*32)];
	assign S1i[1151-((36-30)*32) : 1152-((36-15)*32)] = S0ix[1151-((36-30)*32) : 1152-((36-15)*32)];

	assign S2i[1152-((36-30)*32) +: 32] = S2[127:96];
	assign S2i[1152-((36-31)*32) +: 32] = S2[95:64];
	assign S2i[1152-((36-32)*32) +: 32] = S2[63:32];
	assign S2i[1152-((36-33)*32) +: 32] = S2[31:0];
	assign S2i[1152-((36-27)*32) +: 32] = S1ix[1152-((36-27)*32) +: 32] ^ S2[95:64];
	assign S2i[1152-((36-28)*32) +: 32] = S1ix[1152-((36-28)*32) +: 32] ^ S2[63:32];
	assign S2i[1152-((36-29)*32) +: 32] = S1ix[1152-((36-29)*32) +: 32] ^ S2[31:0];
	assign S2i[1152-((36- 9)*32) +: 32] = S1ix[1152-((36- 9)*32) +: 32] ^ S2[95:64];
	assign S2i[1152-((36-10)*32) +: 32] = S1ix[1152-((36-10)*32) +: 32] ^ S2[63:32];
	assign S2i[1152-((36-11)*32) +: 32] = S1ix[1152-((36-11)*32) +: 32] ^ S2[31:0];
	assign S2i[1151-((36- 9)*32) : 1152-((36-0)*32)] = S1ix[1151-((36- 9)*32) : 1152-((36-0)*32)];
	assign S2i[1151-((36-27)*32) : 1152-((36-12)*32)] = S1ix[1151-((36-27)*32) : 1152-((36-12)*32)];
	assign S2i[1151-((36-36)*32) : 1152-((36-34)*32)] = S1ix[1151-((36-36)*32) : 1152-((36-34)*32)];

	assign S3i[1152-((36-27)*32) +: 32] = S3[127:96];
	assign S3i[1152-((36-28)*32) +: 32] = S3[95:64];
	assign S3i[1152-((36-29)*32) +: 32] = S3[63:32];
	assign S3i[1152-((36-30)*32) +: 32] = S3[31:0];
	assign S3i[1152-((36-24)*32) +: 32] = S2ix[1152-((36-24)*32) +: 32] ^ S3[95:64];
	assign S3i[1152-((36-25)*32) +: 32] = S2ix[1152-((36-25)*32) +: 32] ^ S3[63:32];
	assign S3i[1152-((36-26)*32) +: 32] = S2ix[1152-((36-26)*32) +: 32] ^ S3[31:0];
	assign S3i[1152-((36- 6)*32) +: 32] = S2ix[1152-((36- 6)*32) +: 32] ^ S3[95:64];
	assign S3i[1152-((36- 7)*32) +: 32] = S2ix[1152-((36- 7)*32) +: 32] ^ S3[63:32];
	assign S3i[1152-((36- 8)*32) +: 32] = S2ix[1152-((36- 8)*32) +: 32] ^ S3[31:0];
	assign S3i[1151-((36- 6)*32) : 1152-((36-0)*32)] = S2ix[1151-((36- 6)*32) : 1152-((36-0)*32)];
	assign S3i[1151-((36-24)*32) : 1152-((36-9)*32)] = S2ix[1151-((36-24)*32) : 1152-((36-9)*32)];
	assign S3i[1151-((36-36)*32) : 1152-((36-31)*32)] = S2ix[1151-((36-36)*32) : 1152-((36-31)*32)];

	assign S4i[1152-((36-24)*32) +: 32] = S4[127:96];
	assign S4i[1152-((36-25)*32) +: 32] = S4[95:64];
	assign S4i[1152-((36-26)*32) +: 32] = S4[63:32];
	assign S4i[1152-((36-27)*32) +: 32] = S4[31:0];
	assign S4i[1151-((36-24)*32) : 1152-((36-0)*32)] = S3ix[1151-((36-24)*32) : 1152-((36-0)*32)];
	assign S4i[1151-((36-36)*32) : 1152-((36-28)*32)] = S3ix[1151-((36-36)*32) : 1152-((36-28)*32)];

	smix smix0(clk, S0i[1152-((36-33)*32) +: 32], S0i[1152-((36-34)*32) +: 32], S0i[1152-((36-35)*32) +: 32], S0i[1152-((36- 0)*32) +: 32], S1);
	smix smix1(clk, S1i[1152-((36-30)*32) +: 32], S1i[1152-((36-31)*32) +: 32], S1i[1152-((36-32)*32) +: 32], S1i[1152-((36-33)*32) +: 32], S2);
	smix smix2(clk, S2i[1152-((36-27)*32) +: 32], S2i[1152-((36-28)*32) +: 32], S2i[1152-((36-29)*32) +: 32], S2i[1152-((36-30)*32) +: 32], S3);
	smix smix3(clk, S3i[1152-((36-24)*32) +: 32], S3i[1152-((36-25)*32) +: 32], S3i[1152-((36-26)*32) +: 32], S3i[1152-((36-27)*32) +: 32], S4);

	assign O = { S4i[767:0], S4i[1151:768] };
	
	always @ (posedge clk) begin
		
		S0ixx <= S0i;
		S1ixx <= S1i;
		S2ixx <= S2i;
		S3ixx <= S3i;

		S0ix <= S0ixx;
		S1ix <= S1ixx;
		S2ix <= S2ixx;
		S3ix <= S3ixx;

	end

endmodule

module close_1 (
	input clk,
	input [1151:0] S,
	output [1151:0] out
);

	wire [127:0] S1;
	wire [1151:0] S0i, O;
	reg [1151:0] S0ix;
	reg [1151:0] S0ixx;

	assign S0i[1152-((36- 0)*32) +: 32] = S[1152-((36- 0)*32) +: 32] ^ S[1152-((36- 4)*32) +: 32];
	assign S0i[1152-((36- 1)*32) +: 32] = S[1152-((36- 1)*32) +: 32] ^ S[1152-((36- 5)*32) +: 32];
	assign S0i[1152-((36- 2)*32) +: 32] = S[1152-((36- 2)*32) +: 32] ^ S[1152-((36- 6)*32) +: 32];
	assign S0i[1152-((36-18)*32) +: 32] = S[1152-((36-18)*32) +: 32] ^ S[1152-((36- 4)*32) +: 32];
	assign S0i[1152-((36-19)*32) +: 32] = S[1152-((36-19)*32) +: 32] ^ S[1152-((36- 5)*32) +: 32];
	assign S0i[1152-((36-20)*32) +: 32] = S[1152-((36-20)*32) +: 32] ^ S[1152-((36- 6)*32) +: 32];
	assign S0i[1151-((36-18)*32) : 1152-((36-3)*32)] = S[1151-((36-18)*32) : 1152-((36-3)*32)];
	assign S0i[1151-((36-36)*32) : 1152-((36-21)*32)] = S[1151-((36-36)*32) : 1152-((36-21)*32)];

	smix smix0(clk, S0i[1152-((36-0)*32) +: 32], S0i[1152-((36-1)*32) +: 32], S0i[1152-((36-2)*32) +: 32], S0i[1152-((36-3)*32) +: 32], S1);
	
	assign O = { S0ix[1151:128], S1[31:0], S1[63:32], S1[95:64], S1[127:96] };
	assign out = { O[1055:0], O[1151:1056] };
	
	always @ (posedge clk) begin
		
		S0ixx <= S0i;
		S0ix <= S0ixx;

	end

endmodule

module close_2 (
	input clk,
	input [1151:0] S,
	output [1151:0] O
);

	wire [127:0] S1, S2, S3, S4;

	wire [1151:0] S0i,S1i,S2i,S3i,S4i;
	reg [1151:0] S0ix,S1ix,S2ix,S3ix;
	reg [1151:0] S0ixx,S1ixx,S2ixx,S3ixx;

	assign S0i[1152-((36-13)*32) +: 32] = S[1152-((36- 4)*32) +: 32] ^ S[1152-((36- 0)*32) +: 32];
	assign S0i[1152-((36-18)*32) +: 32] = S[1152-((36- 9)*32) +: 32] ^ S[1152-((36- 0)*32) +: 32];
	assign S0i[1152-((36-27)*32) +: 32] = S[1152-((36-18)*32) +: 32] ^ S[1152-((36- 0)*32) +: 32];
	assign S0i[1152-((36- 0)*32) +: 32] = S[1152-((36-27)*32) +: 32] ^ S[1152-((36- 0)*32) +: 32];
	assign S0i[1151-((36- 9)*32) : 1152-((36- 1)*32)] = S[1151-((36-36)*32) : 1152-((36-28)*32)];
	assign S0i[1151-((36-13)*32) : 1152-((36- 9)*32)] = S[1151-((36- 4)*32) : 1152-((36- 0)*32)];
	assign S0i[1151-((36-18)*32) : 1152-((36-14)*32)] = S[1151-((36- 9)*32) : 1152-((36- 5)*32)];
	assign S0i[1151-((36-27)*32) : 1152-((36-19)*32)] = S[1151-((36-18)*32) : 1152-((36-10)*32)];
	assign S0i[1151-((36-36)*32) : 1152-((36-28)*32)] = S[1151-((36-27)*32) : 1152-((36-19)*32)];

	assign S1i[1152-((36- 9)*32) +: 32] = S1[127:96];
	assign S1i[1152-((36-10)*32) +: 32] = S1[95:64];
	assign S1i[1152-((36-11)*32) +: 32] = S1[63:32];
	assign S1i[1152-((36-12)*32) +: 32] = S1[31:0];
	assign S1i[1152-((36-13)*32) +: 32] = S0ix[1152-((36- 4)*32) +: 32] ^ S1[127:96];
	assign S1i[1152-((36-19)*32) +: 32] = S0ix[1152-((36-10)*32) +: 32] ^ S1[127:96];
	assign S1i[1152-((36-27)*32) +: 32] = S0ix[1152-((36-18)*32) +: 32] ^ S1[127:96];
	assign S1i[1152-((36- 0)*32) +: 32] = S0ix[1152-((36-27)*32) +: 32] ^ S1[127:96];
	assign S1i[1151-((36- 9)*32) : 1152-((36- 1)*32)] = S0ix[1151-((36-36)*32) : 1152-((36-28)*32)];
	assign S1i[1151-((36-19)*32) : 1152-((36-14)*32)] = S0ix[1151-((36-10)*32) : 1152-((36- 5)*32)];
	assign S1i[1151-((36-27)*32) : 1152-((36-20)*32)] = S0ix[1151-((36-18)*32) : 1152-((36-11)*32)];
	assign S1i[1151-((36-36)*32) : 1152-((36-28)*32)] = S0ix[1151-((36-27)*32) : 1152-((36-19)*32)];

	assign S2i[1152-((36- 9)*32) +: 32] = S2[127:96];
	assign S2i[1152-((36-10)*32) +: 32] = S2[95:64];
	assign S2i[1152-((36-11)*32) +: 32] = S2[63:32];
	assign S2i[1152-((36-12)*32) +: 32] = S2[31:0];
	assign S2i[1152-((36-13)*32) +: 32] = S1ix[1152-((36- 4)*32) +: 32] ^ S2[127:96];
	assign S2i[1152-((36-19)*32) +: 32] = S1ix[1152-((36-10)*32) +: 32] ^ S2[127:96];
	assign S2i[1152-((36-28)*32) +: 32] = S1ix[1152-((36-19)*32) +: 32] ^ S2[127:96];
	assign S2i[1152-((36- 0)*32) +: 32] = S1ix[1152-((36-27)*32) +: 32] ^ S2[127:96];
	assign S2i[1151-((36- 9)*32) : 1152-((36- 1)*32)] = S1ix[1151-((36-36)*32) : 1152-((36-28)*32)];
	assign S2i[1151-((36-19)*32) : 1152-((36-14)*32)] = S1ix[1151-((36-10)*32) : 1152-((36- 5)*32)];
	assign S2i[1151-((36-28)*32) : 1152-((36-20)*32)] = S1ix[1151-((36-19)*32) : 1152-((36-11)*32)];
	assign S2i[1151-((36-36)*32) : 1152-((36-29)*32)] = S1ix[1151-((36-27)*32) : 1152-((36-20)*32)];

	assign S3i[1152-((36- 9)*32) +: 32] = S3[127:96];
	assign S3i[1152-((36-10)*32) +: 32] = S3[95:64];
	assign S3i[1152-((36-11)*32) +: 32] = S3[63:32];
	assign S3i[1152-((36-12)*32) +: 32] = S3[31:0];
	assign S3i[1152-((36-13)*32) +: 32] = S2ix[1152-((36- 4)*32) +: 32] ^ S3[127:96];
	assign S3i[1152-((36-19)*32) +: 32] = S2ix[1152-((36-10)*32) +: 32] ^ S3[127:96];
	assign S3i[1152-((36-28)*32) +: 32] = S2ix[1152-((36-19)*32) +: 32] ^ S3[127:96];
	assign S3i[1152-((36- 1)*32) +: 32] = S2ix[1152-((36-28)*32) +: 32] ^ S3[127:96];
	assign S3i[1152-((36- 0)*32) +: 32] = S2ix[1152-((36-27)*32) +: 32];
	assign S3i[1151-((36- 9)*32) : 1152-((36- 2)*32)] = S2ix[1151-((36-36)*32) : 1152-((36-29)*32)];
	assign S3i[1151-((36-19)*32) : 1152-((36-14)*32)] = S2ix[1151-((36-10)*32) : 1152-((36- 5)*32)];
	assign S3i[1151-((36-28)*32) : 1152-((36-20)*32)] = S2ix[1151-((36-19)*32) : 1152-((36-11)*32)];
	assign S3i[1151-((36-36)*32) : 1152-((36-29)*32)] = S2ix[1151-((36-27)*32) : 1152-((36-20)*32)];

	assign S4i[1152-((36- 0)*32) +: 32] = S4[127:96];
	assign S4i[1152-((36- 1)*32) +: 32] = S4[95:64];
	assign S4i[1152-((36- 2)*32) +: 32] = S4[63:32];
	assign S4i[1152-((36- 3)*32) +: 32] = S4[31:0];
	assign S4i[1151-((36-36)*32) : 1152-((36- 4)*32)] = S3ix[1151-((36-36)*32) : 1152-((36- 4)*32)];
	
	smix smix0 (clk, S0i[1152-((36-0)*32) +: 32], S0i[1152-((36-1)*32) +: 32], S0i[1152-((36-2)*32) +: 32], S0i[1152-((36-3)*32) +: 32], S1);
	smix smix1 (clk, S1i[1152-((36-0)*32) +: 32], S1i[1152-((36-1)*32) +: 32], S1i[1152-((36-2)*32) +: 32], S1i[1152-((36-3)*32) +: 32], S2);
	smix smix2 (clk, S2i[1152-((36-0)*32) +: 32], S2i[1152-((36-1)*32) +: 32], S2i[1152-((36-2)*32) +: 32], S2i[1152-((36-3)*32) +: 32], S3);
	smix smix3 (clk, S3i[1152-((36-1)*32) +: 32], S3i[1152-((36-2)*32) +: 32], S3i[1152-((36-3)*32) +: 32], S3i[1152-((36-4)*32) +: 32], S4);
	
	assign O = S4i;
	
	always @ (posedge clk) begin

		S0ixx <= S0i;
		S1ixx <= S1i;
		S2ixx <= S2i;
		S3ixx <= { S3i[31:0], S3i[1151:32] };

		S0ix <= S0ixx;
		S1ix <= S1ixx;
		S2ix <= S2ixx;
		S3ix <= S3ixx;

	end

endmodule
